1 ! 1412
2 " 1344
3 $ 2
4 % 5
5 & 5
6 ' 19
7 ( 889
8 ) 953
9 ): 47
10 + 5
11 , 19817
12 - 1778
13 -(EN 1
14 -(ES 1
15 -54 1
16 -En 1
17 -bearbetning 1
18 -er 1
19 -företag 1
20 -kravet 1
21 -organ 3
22 -politik 1
23 -resurserna 1
24 -är 1
25 . 22037
26 .. 1
27 ... 108
28 .... 1
29 .adp 1
30 .lpk 1
31 .mdb 1
32 .odc 1
33 .udl 1
34 .xml 1
35 .xsd 1
36 .xsl-fil 2
37 / 68
38 0 1
39 0,01 3
40 0,4 1
41 0,6 1
42 0,7 4
43 00.05 1
44 000 102
45 000-3 1
46 008 2
47 0113 1
48 0550 1
49 0652 1
50 09.00 1
51 1 115
52 1,2 2
53 1,27 1
54 1,4 1
55 1,5 1
56 1,7 2
57 1,8 1
58 1,84 1
59 1,9 1
60 1-2 1
61 1-3 1
62 1-bil 1
63 1-fonderna 1
64 1-land 1
65 1-område 1
66 1-områden 1
67 1-områdena 3
68 1-området 1
69 1-region 1
70 1-regioner 2
71 1-regionerna 3
72 1-status 2
73 1-stöden 1
74 1/3 1
75 10 48
76 10,9 1
77 10.000 1
78 10.40 1
79 100 25
80 100-procentig 1
81 101 1
82 102 2
83 103 2
84 104 2
85 105 4
86 106 1
87 107 3
88 107:e 1
89 108 2
90 11 33
91 11,3 1
92 11.00 11
93 11.1 3
94 11.10 1
95 11.25 1
96 11.30 7
97 110 2
98 110:e 1
99 11195/1/1999 1
100 112 1
101 11287/1/1999 1
102 112:e 1
103 114 1
104 115 1
105 116:e 1
106 119:e 1
107 11d 1
108 12 34
109 12.00 27
110 12.25 1
111 12.30 1
112 12.40 1
113 12/99 3
114 120 2
115 122 1
116 123 2
117 1244 6
118 12485/1/1999 1
119 12487/1/1999 1
120 125 1
121 1257/99 1
122 1260 1
123 1260/1999om 1
124 1260/99 1
125 127 1
126 1284 2
127 129 1
128 13 52
129 13,5 2
130 13,9 1
131 13-14 3
132 13.05 1
133 13.23 1
134 13.40 1
135 13.55 1
136 130 2
137 133.2 1
138 137 1
139 138 1
140 138.4 1
141 14 45
142 14,7 1
143 14.10 1
144 140 2
145 1408 1
146 14094/1999 2
147 142 1
148 143 1
149 1448 1
150 15 50
151 15,2 1
152 15,4 1
153 15.00 5
154 15.45 1
155 15.50 1
156 150 7
157 152 11
158 158 5
159 158.1 1
160 159 1
161 16 27
162 16.05 1
163 16.30 2
164 1626 1
165 1626/94 1
166 1638 1
167 164 2
168 166 2
169 167 3
170 17 18
171 17.30 1
172 170 1
173 174 1
174 1762 2
175 177 2
176 1775 1
177 178 1
178 18 29
179 18.00 4
180 180 1
181 1800-talet 2
182 1809 2
183 19 10
184 19.05 1
185 19.15 1
186 19.30 1
187 19.40 1
188 19.50 1
189 190 2
190 1900 1
191 1900-talet 4
192 191 1
193 1910 3
194 1917 1
195 1923 1
196 1929 3
197 193 1
198 1930-talet 2
199 194 1
200 1945 1
201 1947 3
202 1948 1
203 1949 2
204 195 1
205 1952 1
206 1953 1
207 1955 1
208 1957 6
209 1958 1
210 1959 1
211 1960 2
212 1967 7
213 1969 2
214 1970 1
215 1973 1
216 1974 3
217 1975 2
218 1976 1
219 1977 2
220 1978 1
221 1979 2
222 1980-talet 2
223 1981 1
224 1982 2
225 1983 1
226 1984 4
227 1986 7
228 1987 3
229 1988 4
230 1989 6
231 1990 12
232 1990-talet 6
233 1991 5
234 1992 15
235 1993 16
236 1993-1995 2
237 1994 20
238 1994-1999 5
239 1995 24
240 1995-1997 1
241 1996 28
242 1996-1997 1
243 1997 56
244 1997/0067(COD 2
245 1997/0194(COD 2
246 1997/0352(CNS 1
247 1997/0370(COD 2
248 1997/0371(COD 2
249 1998 57
250 1998-2002 2
251 1998/0097(COD 1
252 1998/0106(COD 2
253 1998/0141 2
254 1998/0169(COD 2
255 1998/0242(COD 1
256 1998/0249(COD 1
257 1998/0324(COD 2
258 1999 154
259 1999-2000 1
260 1999-2004 1
261 1999-2006 1
262 1999/0012(COD 1
263 1999/0013(CNS 1
264 1999/0015(COD 1
265 1999/0020(COD 1
266 1999/0083 1
267 1999/0090(COD 1
268 1999/0168(CNS 2
269 1999/0196(CNS 2
270 1999/0199(CNS 2
271 1999/0218(CNS 1
272 1999/0222(CNS 1
273 1999/0224(CNS 1
274 1999/0228(CNS 1
275 1999/0240(CNS 2
276 1999/0803(CNS 1
277 1999/0805(CNS 1
278 1999/0806(CNS 1
279 1999/0809(CNS 1
280 1999/0821(CNS 2
281 1999/0825(CNS 2
282 1999/2115(COS 1
283 1999/2121(COS 2
284 1999/2123(COS 1
285 1999/2127(COS 1
286 1999/2150(COS 2
287 1999/2155(COS 2
288 1999/2182(COS 2
289 1999/2186(COS 1
290 1999/468 4
291 2 91
292 2,3 1
293 2,487 1
294 2,5 2
295 2,6 1
296 2,8 3
297 2,9 1
298 2-område 1
299 2-områdena 1
300 2-stöd 1
301 2.1 1
302 2.2 2
303 2.7 2
304 20 54
305 20.15 1
306 20.25 1
307 20.30 2
308 200 16
309 2000 138
310 2000- 1
311 2000-2001 1
312 2000-2004 6
313 2000-2005 8
314 2000-2006 25
315 2000-2010 1
316 2000-buggen 1
317 2000-filformat 3
318 2000-korsetten 1
319 2000-paketet 1
320 2000-platser 1
321 2000-programmet 4
322 2000-talet 5
323 2000-talets 2
324 2000-versionen 1
325 2000/2046(COS 2
326 2001 15
327 2002 35
328 2002- 2
329 2002-filformat 2
330 2003 10
331 2004 4
332 2005 4
333 2006 11
334 2007 2
335 2008 1
336 2010 10
337 2012 3
338 2020 12
339 2025 1
340 2034 1
341 205 1
342 21 16
343 21.00 5
344 21.1 1
345 21.55 1
346 2100 1
347 21:a 5
348 22 19
349 22,5 1
350 22.3 1
351 22.41 1
352 2200 1
353 226 1
354 22a 1
355 23 10
356 23,7 1
357 23-24 2
358 23.50 1
359 23.55 1
360 235- 1
361 24 20
362 24,5 1
363 240 2
364 243 1
365 245 1
366 246 1
367 248 2
368 249 4
369 25 40
370 25,7 1
371 25,9 1
372 25-åriga 1
373 250 3
374 251 1
375 255 4
376 25ºC 1
377 26 17
378 262 1
379 263 1
380 27 11
381 270 3
382 27º 1
383 28 18
384 28,2 1
385 280 4
386 280.4 1
387 28:e 1
388 29 11
389 29,9 2
390 29.4 1
391 299.2 2
392 2l:a 1
393 3 63
394 3,5 1
395 3,604 1
396 3,8 2
397 3,9 1
398 3-4 1
399 3-liter-bilar 1
400 3-liters-bilen 1
401 3.1 1
402 3.8 1
403 3/4 2
404 30 32
405 30,8 1
406 300 11
407 300.3 1
408 3062 1
409 308- 1
410 30:1 1
411 31 21
412 310 1
413 314 1
414 32 10
415 33 10
416 33,4 1
417 332 1
418 34 12
419 34.1.1 1
420 34.2 2
421 340 1
422 344 1
423 347 2
424 35 15
425 35-40 1
426 35-timmarslagen 1
427 35-timmarsvecka 1
428 35-årige 1
429 350 3
430 36 7
431 3605/93 3
432 363 2
433 366 1
434 367 1
435 37 23
436 37.2 5
437 37/60/92 1
438 370 3
439 378 2
440 38 12
441 388 2
442 39 10
443 394/2000 1
444 4 72
445 4,3 1
446 4,5 1
447 4,875 1
448 4-5 1
449 4.2 1
450 4.5 1
451 40 31
452 40-aktien 1
453 40-procentigt 1
454 400 12
455 41 8
456 410 1
457 42 8
458 42.2 1
459 42.5 1
460 43 12
461 43- 1
462 44 10
463 444 2
464 45 20
465 45-varvare 1
466 451 1
467 453 1
468 46 6
469 462 1
470 47 7
471 476 1
472 47e 1
473 48 9
474 49 8
475 4:ans 1
476 5 57
477 5,1 1
478 5,2 1
479 5,3 1
480 5,35 1
481 5,5 2
482 5,8 1
483 5-10 1
484 5.4 1
485 50 44
486 50- 1
487 50-tal 1
488 50-talskulturen 1
489 50-årsdagen 1
490 50-årsjubileum 1
491 50-årsjubiléum 1
492 500 12
493 5060/1999 1
494 51 3
495 5116/1999 2
496 519 1
497 52 3
498 520 2
499 522 1
500 53 6
501 535 2
502 54 4
503 540 1
504 541 1
505 55 5
506 551 1
507 552 1
508 55:e 2
509 55º 1
510 56 5
511 56:e 3
512 57 2
513 57,5 1
514 5713/1999 1
515 58 2
516 59 4
517 5b 3
518 5b-området 1
519 6 64
520 6,07 1
521 6,4 2
522 6.1 4
523 60 21
524 60-talet 1
525 600 4
526 60:1 1
527 60º 1
528 61 1
529 613 8
530 615 1
531 62 3
532 623 2
533 63 2
534 64 1
535 65 3
536 650 1
537 6500 1
538 658 1
539 66 1
540 66,3 1
541 67 3
542 68 2
543 685/95 1
544 69 2
545 69.2 2
546 7 73
547 7,2 2
548 7,42 1
549 7,5 1
550 7-9 1
551 7.1 3
552 7.2 1
553 70 10
554 70/524 7
555 700 10
556 70:e 1
557 71 8
558 717 1
559 72 2
560 72:a 2
561 73 2
562 73,9 1
563 74 1
564 747:an 1
565 74:1 1
566 75 11
567 76 4
568 768 1
569 77 3
570 78 2
571 784 1
572 79 4
573 79/409 1
574 8 38
575 80 30
576 80-90 1
577 80-procentiga 1
578 80-talet 1
579 800 8
580 8095/1/1999 2
581 81 7
582 81(rev 1
583 81.1 5
584 81.3 5
585 82 8
586 83 3
587 830 1
588 84 2
589 85 9
590 85/611 4
591 850 9
592 850/98 1
593 86 4
594 87 5
595 87.1 1
596 87.2 1
597 88 4
598 88/591 2
599 89 3
600 9 35
601 9,2 1
602 9,5 2
603 9.00 1
604 9.1 1
605 90 17
606 90-talet 2
607 90/220 6
608 90/424 3
609 900 3
610 9085/3/1999 2
611 91 2
612 91/68 2
613 9178/1999 1
614 919 1
615 92 1
616 92/43 1
617 93 2
618 93/53 2
619 93/75 1
620 94 5
621 94/55 2
622 94/728 1
623 95 21
624 95/35 1
625 96 1
626 96/23 1
627 96/35 3
628 96/71 2
629 96/96 1
630 9614/1999 1
631 9636/1999 1
632 97 2
633 97-filformat 1
634 97/67 1
635 97/99 1
636 9767 1
637 97:e 1
638 98 3
639 99 2
640 : 1022
641 ; 381
642 ? 948
643 A 13
644 A-tjänstemän 1
645 A. 2
646 A32 1
647 A4-0029/2000 1
648 A4-0072/97 1
649 A5-0001/2000 1
650 A5-0002/2000 1
651 A5-0003/2000 2
652 A5-0004/2000 1
653 A5-0006/00 1
654 A5-0006/2000 2
655 A5-0007/2000 3
656 A5-0008/2000 3
657 A5-0009/2000 2
658 A5-0010/2000 2
659 A5-0011/2000 2
660 A5-0012/2000 2
661 A5-0013/2000 2
662 A5-0014/2000 2
663 A5-0015/2000 2
664 A5-0015/2000)av 1
665 A5-0016/2000 2
666 A5-0017/2000 3
667 A5-0018/2000 2
668 A5-0019/2000 3
669 A5-0020/2000 3
670 A5-0021/2000 2
671 A5-0022/2000 2
672 A5-0023/2000 3
673 A5-0025/2000 2
674 A5-0026/2000 1
675 A5-0027/2000 3
676 A5-0028/2000 1
677 A5-0029/2000 2
678 A5-0031/2000 3
679 A5-0032/2000 3
680 A5-0033/2000 3
681 A5-0034/2000 3
682 A5-0035/2000 1
683 A5-0036/2000 2
684 A5-0037/2000 1
685 A5-0038/2000 2
686 A5-0039/2000 1
687 A5-0040/2000 1
688 A5-0041/2000 2
689 A5-0043/2000 2
690 A5-0048/2000 1
691 A5-0051/2000 1
692 A5-0069/1999 1
693 A5-0073/1999 1
694 A5-0078/1999 1
695 A5-0087/1999 1
696 A5-0104/1999 2
697 A5-0105/1999 2
698 A5-0106/1999 1
699 A5-0107/1999 2
700 A5-0108/1999 2
701 A5­0030/2000 1
702 ABB 4
703 ABB-Alsthom 2
704 ABB-Alstom 2
705 ABC 1
706 ADOX 1
707 ADR 1
708 AKTUELLA 2
709 ALE 1
710 ALE- 1
711 ALE-gruppen 2
712 ANSI 16
713 ANSI-89 10
714 ANSI-92 11
715 ANSI-92-frågor 1
716 ANSI-92-läge 1
717 ANSI-syntax 1
718 AVC 2
719 AVS 7
720 AVS-EU 3
721 AVS-EU-avtalet 1
722 AVS-EU-partnerskapet 1
723 AVS-EU:s 11
724 AVS-grannar 1
725 AVS-gruppen 1
726 AVS-gruppens 1
727 AVS-land 1
728 AVS-landet 1
729 AVS-länder 5
730 AVS-länderna 35
731 AVS-ländernas 9
732 AVS-partner 3
733 AVS-samarbetet 3
734 AVS-staterna 3
735 AVS-staternas 2
736 Absaloms 1
737 Absolut 3
738 Accepterandet 1
739 Access 32
740 Access-databas 5
741 Access-databaser 2
742 Access-databasobjekt 1
743 Access-fil 2
744 Access-filen 1
745 Access-filer 1
746 Access-projekt 3
747 Act 2
748 Action 1
749 Adam 1
750 Adamson 7
751 Adana 1
752 Adapt 2
753 Adapt- 1
754 Adapt-projekt 1
755 Additionalitet 1
756 Adelaide 1
757 Adenauer 1
758 Adjö 1
759 Administration 1
760 Admiral 1
761 Adolf 2
762 Adriatiska 3
763 Advanced 1
764 Advertising 1
765 Advokaten 1
766 Afrika 53
767 Afrikanska 2
768 Afrikas 2
769 Afrodites 1
770 Agenda 20
771 Agents 1
772 Agliettas 1
773 Agrifin-rådet 1
774 Agustaaffären 1
775 Aha 1
776 Ahern 8
777 Ahmed 1
778 Aids 1
779 Aidsbehandlingar 1
780 Aidsproblemet 1
781 Air 2
782 Aires 1
783 Airways 1
784 Akkuyu 2
785 Akköy 1
786 Aktiviteterna 1
787 Alan 1
788 Alavanos 9
789 Albacète 1
790 Albaner 1
791 Albanien 13
792 Albert 1
793 Albright 1
794 Aldrig 5
795 Alex 3
796 Alexander 3
797 Alexandra 2
798 Alexandros 1
799 Alfanjurt 1
800 Alfen 1
801 Algarve 1
802 Algeriet 1
803 Algeriets 1
804 Algonquin 3
805 Alicante 2
806 Alicante-byrån 1
807 Alice 3
808 Alkartasuna 1
809 Alkoholmonopol 1
810 Alkoholpolitiken 1
811 All 4
812 Alla 84
813 Alldeles 6
814 Allen 1
815 Allesammans 1
816 Allmänheten 2
817 Allmänna 1
818 Allmänt 3
819 Allra 1
820 Allt 44
821 Alltför 3
822 Alltid 1
823 Allting 3
824 Alltsedan 3
825 Alltså 5
826 Almería 4
827 Alonso 1
828 Alperna 1
829 Alsace 4
830 Alsthom 1
831 Alstom 2
832 Altener 8
833 Altener-program 1
834 Altener-programmet 9
835 Alternativet 1
836 Alyssandrakis 3
837 Amadeus 1
838 Amado 4
839 Ambitionen 1
840 Ambrogio 1
841 Amerika 5
842 Amerikanerna 1
843 Amerikas 5
844 Amiens 1
845 Amins 1
846 Ammokosto 1
847 Amnesty 1
848 Amoco 2
849 Amoco-Cádiz 1
850 Amoko 5
851 Amos 1
852 Amsterdam 17
853 Amsterdamfördrag 1
854 Amsterdamfördraget 46
855 Amsterdamfördragets 1
856 Amsterdamresterna 1
857 Amsterdams 1
858 Andalusien 14
859 Andelen 1
860 Andersens 1
861 Andersonbetänkandet 1
862 Andersson 19
863 Anderssonbetänkandet 3
864 Anderssons 8
865 Andliga 1
866 Andra 16
867 Andrabehandlingsrekommendation 5
868 Andrej 14
869 Andrew 2
870 Angelilli 1
871 Angola 33
872 Angolafrågan 1
873 Angolas 2
874 Angående 57
875 Anhållandena 1
876 Ankara 5
877 Ankaras 1
878 Anledningen 2
879 Anläggning 1
880 Anmälningsplikten 1
881 Anna 1
882 Annan 1
883 Annars 9
884 Anpassa 2
885 Anpassningen 1
886 Anser 14
887 Anslagen 1
888 Anslagsbeloppet 1
889 Ansträngningarna 1
890 Anställda 1
891 Ansvaret 4
892 Ansvariga 1
893 Ansvarsfrihet 1
894 Ansvarsfriheten 1
895 Antagandet 1
896 Antal 2
897 Antalet 3
898 Antar 1
899 Antas 1
900 Antibiotika 1
901 Antingen 6
902 Antwerpen 1
903 António 3
904 Anvers 1
905 Använda 5
906 Användandet 1
907 Användare 3
908 Användaren 3
909 Användarna 2
910 Användning 1
911 Användningen 4
912 Aparicio 1
913 Apollo 1
914 Apostrofen 1
915 Applications 1
916 Applåder 17
917 Apropå 3
918 Arabic 1
919 Arabrepubliken 1
920 Arabvärldens 1
921 Arafat 1
922 Arafats 1
923 Arbete 1
924 Arbetet 5
925 Arbetskultur 1
926 Arbetslöshet 1
927 Arbetslösheten 2
928 Arbetslöshetssiffrorna 1
929 Arbetsmarknad 1
930 Arbetsmarknaden 1
931 Arbetsmarknadsministeriet 1
932 Arbetspasset 1
933 Arbetsplan 2
934 Arbetsplanen 1
935 Arbetstagarna 1
936 Arbetstidsdirektivet 1
937 Arbetsvillkoren 1
938 Argumentet 1
939 Ari 1
940 Ariane 3
941 Arizona 5
942 Arkimedes 1
943 Arkiv-menyn 1
944 Armarna 1
945 Armenien 14
946 Arms 1
947 Arousa 1
948 Artas 1
949 Arthur 1
950 Artikel 6
951 Artikeln 1
952 Artiklarna 2
953 Arts 1
954 Asahe 2
955 Asien 4
956 Aspe-dalen 1
957 Aspects 1
958 Assad 2
959 Associations 2
960 Asturien 1
961 Ataturk-dammarna 1
962 Atatürkdammarna 1
963 Aten 1
964 Athen 1
965 Athena 4
966 Atlantalliansen 1
967 Atlantbågens 1
968 Atlanten 13
969 Atlantic 1
970 Atlantkust 1
971 Atlantkusten 3
972 Atlantkustens 1
973 Att 117
974 Attacken 1
975 Attwool 3
976 Attwooll 6
977 Attwoolls 1
978 Atxalandabaso 2
979 Aubert 1
980 Auerbach 2
981 Aung 1
982 Auroi 2
983 Auschwitz 2
984 Auster 22
985 Austers 7
986 Australien 1
987 Authoring 1
988 Auto 1
989 Autofilter 1
990 Autofiltrering 1
991 Auvergne 1
992 Av 75
993 Avbrottet 1
994 Avbrytande 3
995 Avenue 3
996 Avfallet 1
997 Avgången 1
998 Aviano 1
999 Avlägset 1
1000 Avreglering 2
1001 Avregleringen 2
1002 Avsaknaden 1
1003 Avsatta 1
1004 Avser 1
1005 Avsevärda 1
1006 Avsikten 3
1007 Avskaffandet 1
1008 Avslutande 1
1009 Avslutningsvis 41
1010 Avslöja 1
1011 Avtal 1
1012 Avtalen 1
1013 Avtalens 1
1014 Avtalet 9
1015 Azerbajdzjan 1
1016 Aziz 1
1017 Aznar 5
1018 Azorerna 5
1019 B 9
1020 B. 4
1021 B1-382 1
1022 B1-500 1
1023 B2-5122 1
1024 B5-0003/2000 2
1025 B5-0009/2000 2
1026 B5-0010/2000 1
1027 B5-0011/2000 1
1028 B5-0012/2000 1
1029 B5-0040/99 1
1030 B5-0041/99 1
1031 B5-0125/2000 1
1032 B5-0132/2000 1
1033 B5-0136/2000 1
1034 B5-0140/2000 1
1035 B5-0141/2000 1
1036 B5-0142/2000 1
1037 B5-0148/2000 1
1038 B5-0149/2000 1
1039 B5-0150/2000 1
1040 B5-0151/2000 1
1041 B5-0152/2000 1
1042 B5-0153/2000 1
1043 B5-0154/2000 1
1044 B5-0155/2000 1
1045 B5-0156/2000 1
1046 B5-0157/2000 1
1047 B5-0158/2000 1
1048 B5-0159/2000 1
1049 B5-0160/2000 1
1050 B5-0161/2000 1
1051 B5-0162/2000 1
1052 B5-0163/2000 1
1053 B5-0164/2000 1
1054 B5-0165/2000 1
1055 B5-0166/2000 1
1056 B5-0167/2000 1
1057 B5-0168/2000 1
1058 B5-0169/2000 1
1059 B5-0170/2000 1
1060 B5-0171/2000 1
1061 B5-0172/2000 1
1062 B5-0173/2000 1
1063 B5-0174/2000 1
1064 B5-0175/2000 1
1065 B5-0176/2000 1
1066 B5-0177/2000 1
1067 B5-0178/2000 1
1068 B5-0179/2000 1
1069 B5-0180/2000 1
1070 B5-0181/2000 2
1071 B7 1
1072 B7-0 1
1073 B7-04 1
1074 B7-4011 1
1075 B7-4012 1
1076 B7-6201 1
1077 BAT 1
1078 BBC 4
1079 BBC-intervju 1
1080 BBC:s 1
1081 BNI 13
1082 BNI-tillväxt 1
1083 BNP 9
1084 BP 1
1085 BRAY 1
1086 BRÅDSKANDE 2
1087 BSE 13
1088 BSE-epidemin 1
1089 BSE-krisen 4
1090 BSE-tester 1
1091 BSE-typ 1
1092 BSE-utskott 1
1093 BSE-utskottets 1
1094 Babitskij 15
1095 Babitskijaffären 1
1096 Babitskijs 3
1097 Baconsmörgåsarna 1
1098 Bakom 7
1099 Balfe 1
1100 Balford-förklaringen 1
1101 Balkan 51
1102 Balkanhalvöns 1
1103 Balkanländerna 2
1104 Balkanregionen 1
1105 Balkanrepublik 1
1106 Balkans 4
1107 Banantvisten 1
1108 Bandet 1
1109 Bangemann 1
1110 Bangkok 1
1111 Bank 1
1112 Bankgarantier 1
1113 Bankrutten 1
1114 Banotti 9
1115 Bara 16
1116 Barak 6
1117 Baraks 3
1118 Barcelonaprocess 1
1119 Barcelonaprocessen 1
1120 Barcelonaprocessens 1
1121 Baren 2
1122 Barents 1
1123 Baringdorf 9
1124 Barn 2
1125 Barnet 1
1126 Barnhill 1
1127 Barnier 28
1128 Barniers 4
1129 Barry 1
1130 Bartho 1
1131 Barzanti 1
1132 Barzantibetänkandet 1
1133 Barón 6
1134 Basel 1
1135 Basel-Mulhouse-flygplatsen 1
1136 Basic 2
1137 Basic-projektet 1
1138 Baskien 15
1139 Baskiens 2
1140 Bassam 1
1141 Basse-Normandie 1
1142 Battery 1
1143 Bautista 1
1144 Bay 1
1145 Bayley 4
1146 Bayleys 2
1147 Bazin 1
1148 Beakta 1
1149 Beatles 3
1150 Beazley 1
1151 Bedfordshire 1
1152 Bediener 1
1153 Bedrägeri 1
1154 Bedrägeri- 1
1155 Bedömningen 2
1156 Beets 1
1157 Befolkningarnas 1
1158 Befolkningen 3
1159 Befordringssystemet 1
1160 Begreppet 2
1161 Begränsa 1
1162 Begränsningar 1
1163 Begär 1
1164 Behandlingen 2
1165 Behöver 3
1166 Bekvämlighetsflaggen 2
1167 Bekämpandet 1
1168 Bekämpning 1
1169 Belgien 16
1170 Belgiens 2
1171 Belgrad 8
1172 Belgrads 2
1173 Belize 2
1174 Belzecs 1
1175 Ben-Gurion 3
1176 Benelux 1
1177 Benengeli-kvartetten 1
1178 Berend 9
1179 Berendbetänkandet 1
1180 Berends 2
1181 Berenguer 3
1182 Berg 1
1183 Bergen 6
1184 Berger 11
1185 Bergerbetänkandet 1
1186 Berlin 16
1187 Berlinavtalen 1
1188 Berlinmurens 1
1189 Bern- 1
1190 Bern-konventionen 1
1191 Bernard 12
1192 Bernd 3
1193 Bernie 1
1194 Bernié 1
1195 Beroende 1
1196 Beroendet 1
1197 Beror 1
1198 Berthu 5
1199 Bertinotti 1
1200 Berätta 1
1201 Beskrivningen 1
1202 Beslut 1
1203 Beslutet 9
1204 Beslutsfattandet 1
1205 Besque 1
1206 Bestämmelserna 1
1207 Besättningen 1
1208 Betoningen 1
1209 Beträffande 18
1210 Betty 1
1211 Betydande 1
1212 Betydelsen 1
1213 Betänkande 52
1214 Betänkandena 1
1215 Betänkandet 13
1216 Betänkligheterna 1
1217 Beveridges 1
1218 Beviljandet 1
1219 Beviset 2
1220 Bibel 2
1221 Bibeln 2
1222 Bidraget 1
1223 Big 5
1224 Bilbao 2
1225 Bilder 2
1226 Bilen 1
1227 Bilindustrin 1
1228 Bilkonceptet 1
1229 Bill 1
1230 Billobbyn 2
1231 Biltillverkare 2
1232 Birds 1
1233 Biscaya 1
1234 Biscayabukten 3
1235 Biscayagolfen 4
1236 Biståndet 1
1237 Biståndsgivarens 1
1238 Biståndsnivån 2
1239 Bit 1
1240 Bjerregaard 1
1241 Blak 2
1242 Blanco 3
1243 Bland 14
1244 Blanda 1
1245 Blok 1
1246 Blokland 1
1247 Blooms 1
1248 Blotts 1
1249 Blåfenad 1
1250 Boetticher 1
1251 Bohéme 1
1252 Boken 1
1253 Bokhållaren 1
1254 Bolagsdirektören 1
1255 Bolkestein 19
1256 Bolkesteins 1
1257 Bologna 1
1258 Bom 1
1259 Bomber 1
1260 Bonde 7
1261 Bonino 2
1262 Bonino-listan 1
1263 Booz 1
1264 Bor 1
1265 Borde 8
1266 Bordeaux 1
1267 Borgia 1
1268 Borgin 6
1269 Borgins 2
1270 Borràs 3
1271 Bortanför 1
1272 Bortom 2
1273 Bortre 1
1274 Bortsållning 1
1275 Bos 1
1276 Bosnien 5
1277 Bosnien-Hercegovina 1
1278 Bosnien-Herzegovina 4
1279 Bosniens 1
1280 Bosse 1
1281 Boston 1
1282 Bosättarna 1
1283 Botswana 1
1284 Bourlanges 6
1285 Bouwman 10
1286 Bowe 2
1287 Bowis 2
1288 Boyne 3
1289 Boynes 2
1290 Boynesmynningen 1
1291 Boynesmynningens 1
1292 Bra 1
1293 Braer 2
1294 Braerkatastrofen 1
1295 Brahim 1
1296 Brandenburg 2
1297 Branschen 1
1298 Brasilien 3
1299 Bravery 1
1300 Bray 31
1301 Bremen 1
1302 Brempt 1
1303 Bresjnevs 1
1304 Bretagne 16
1305 Bretagnes 3
1306 Bretonne 1
1307 Brevbäraren 1
1308 Brian 1
1309 Brist 2
1310 Bristen 1
1311 Bristerna 1
1312 British 3
1313 Brittan 1
1314 Brittiska 1
1315 Broadway 3
1316 Broek 1
1317 Brok 18
1318 Brokbetänkandet 2
1319 Broks 4
1320 Bronislav 1
1321 Brottsligheten 1
1322 Brovina 8
1323 Brovinas 1
1324 Brown 1
1325 Brundtland-rapporten 1
1326 Bruno 1
1327 Bryssel 54
1328 Bryssel-I 1
1329 Bryssel-II 1
1330 Brysselartikeln 1
1331 Brysselbyråkrater 1
1332 Brysselbyråkratin 1
1333 Brysselfederalistiskt 1
1334 Brysselfördraget 1
1335 Bryssels 2
1336 Brysselteknokraternas 1
1337 Bränningens 1
1338 Bröderna 1
1339 Budapest 3
1340 Budget- 1
1341 Budgetförordningen 2
1342 Budgetmedlen 1
1343 Budgetplanerna 1
1344 Budgetutskottet 1
1345 Buenos 1
1346 Buesa 5
1347 Bulgarien 8
1348 Bundestag 1
1349 Burkes 2
1350 Burkina 1
1351 Burma 11
1352 Bush 1
1353 Busquin 1
1354 Busquins 2
1355 Bygget 1
1356 Byrne 11
1357 Byrån 7
1358 BÄTTRE 1
1359 Bägge 1
1360 Bästa 1
1361 Bäste 2
1362 Bättre 1
1363 Båda 10
1364 Både 8
1365 Béguin 2
1366 Böcker 1
1367 Böge 6
1368 Böges 2
1369 Böhm 1
1370 Bör 1
1371 Börja 1
1372 Bösch 1
1373 Bülent 2
1374 C 4
1375 C. 4
1376 C4-0018/98 1
1377 C4-0026/1999 2
1378 C4-0212/1999 1
1379 C4-0350/1998 1
1380 C4-0351/1998 1
1381 C4-0352/1999 1
1382 C4-0465/1998 1
1383 C4-0497/98-98/0126 1
1384 C4-0715/98-98/0318(SYN 1
1385 C5-0004/1999 1
1386 C5-0013/2000 1
1387 C5-0014/00 1
1388 C5-0020/1999 1
1389 C5-0040/2000 1
1390 C5-0045/00 1
1391 C5-0045/2000 1
1392 C5-0050/2000 1
1393 C5-0069/1999 1
1394 C5-0081/2000 2
1395 C5-0091/1999 1
1396 C5-0095/1999 1
1397 C5-0112/1999 1
1398 C5-0120/99 1
1399 C5-0122/1999 1
1400 C5-0134/1999 2
1401 C5-0156/1999 2
1402 C5-0166/1999 2
1403 C5-0167/1999 1
1404 C5-0174/1999 2
1405 C5-0176/1999 2
1406 C5-0180/1999 2
1407 C5-0208/1999 2
1408 C5-0209/1999 2
1409 C5-0222/1999 2
1410 C5-0251/99 1
1411 C5-0253/1999 2
1412 C5-0260/1999 1
1413 C5-0302/1999 1
1414 C5-0303/1999 1
1415 C5-0305/1999 1
1416 C5-0308/1999 2
1417 C5-0323/99 1
1418 C5-0327/1999 2
1419 C5-0331/1999 1
1420 C5-0332/1999 2
1421 C5-0333/1999 2
1422 C5-0334/1999 2
1423 C5-0341/1999 2
1424 CAC 3
1425 CECAF:s 1
1426 CEN 8
1427 CEN:s 4
1428 CERN 1
1429 CIA 3
1430 CIP 1
1431 CNS 1
1432 COD 1
1433 COPA 1
1434 CORUS 1
1435 COSV 1
1436 CSS-fil 1
1437 CSU-gruppens 1
1438 CSU:s 2
1439 CTRL-C. 1
1440 CTRL-V. 1
1441 Cadiz 4
1442 Cadiz-katastrofen 2
1443 Cadou 1
1444 Caesarea 1
1445 Caillaux 1
1446 Calais 1
1447 Cambridge 1
1448 Camdessus 1
1449 Campos 1
1450 Camre 1
1451 Camus 1
1452 Canada 1
1453 Candutyp 1
1454 Canyon 3
1455 Canyons 1
1456 Cappuccino 1
1457 Cara-programmet 1
1458 Cardiff 2
1459 Cardiffprocessen 2
1460 Carlo 1
1461 Caroline 1
1462 Casablanca 1
1463 Casaca 1
1464 Casas 2
1465 Cashman 1
1466 Castro-regimen 1
1467 Caudron 1
1468 Cavalese 1
1469 Cederschiöld 13
1470 Cederschiöldbetänkandet 1
1471 Cederschiölds 5
1472 Celsius 3
1473 Cem 1
1474 Central- 11
1475 Centralamerika 2
1476 Centralasiatiska 2
1477 Centralasien 3
1478 Centralasiens 1
1479 Centralbanken 3
1480 Centralbankschefen 1
1481 Centraleuropa 2
1482 Cermis 1
1483 Cervantes 1
1484 Ceyhun 1
1485 Champagne-Ardennes 1
1486 Chanel 1
1487 Change 1
1488 Chapmanfyren 1
1489 Charente 1
1490 Charles 1
1491 Charlie 2
1492 Charlotte 1
1493 Chefen 1
1494 Chevènement 1
1495 Chicago 2
1496 Chile 2
1497 Chiquita 1
1498 Chissano 1
1499 Chris 1
1500 Christine 1
1501 Christopher 4
1502 Church 1
1503 Ciampi-gruppen 1
1504 Circa 1
1505 Cirka 2
1506 Cisterna 6
1507 Clare 1
1508 Claude 3
1509 Clintons 1
1510 Clough 1
1511 Clément 1
1512 Coca 1
1513 Cocilovo 1
1514 Coco 1
1515 Cocoon 1
1516 Coelho 1
1517 Coffee 1
1518 Cohn-Bendit 6
1519 Cola 1
1520 Colombia 2
1521 Comartkommitté 1
1522 Comartkommittén 1
1523 Comité 1
1524 Commission 2
1525 Community 1
1526 Company 1
1527 Companys 1
1528 Compensation 1
1529 Components 5
1530 Components-element 1
1531 Compostela 1
1532 Compson 1
1533 Compsons 1
1534 Conakry 1
1535 Confederation 1
1536 Connaught 1
1537 Connection 1
1538 ConnectionFile 4
1539 ConnectionString 6
1540 Consortium 1
1541 Constabulary 1
1542 Contre 1
1543 Copeland 3
1544 Copyright 1
1545 Corbett 7
1546 Core-projektet 1
1547 Corinne 1
1548 Cork 3
1549 Cornelissen 1
1550 Cornwall 1
1551 Corporate 1
1552 Corpus 1
1553 Corrie 17
1554 Corrie-betänkandet 1
1555 Corriebetänkandet 1
1556 Corriebetänkandets 1
1557 Cossutta 1
1558 Costa 11
1559 Council 1
1560 Cox 8
1561 Coûteaux 1
1562 Crab 1
1563 Crespo 2
1564 Crespos 2
1565 Cresson 2
1566 Crisex 1
1567 Crowley 3
1568 Cummings 3
1569 Cunard 2
1570 Cunardbolaget 1
1571 Cunards 1
1572 Cunha 1
1573 Cunhabetänkandet 1
1574 Cunhas 1
1575 Curie-stipendier 1
1576 Curtis 2
1577 Cushnahan 1
1578 Cusí 1
1579 Cusís 2
1580 Cuxhaven 1
1581 Cyaniden 1
1582 Cymru 1
1583 Cypern 73
1584 Cypernfrågan 6
1585 Cypernkonflikten 1
1586 Cypernproblemet 1
1587 Cyperns 14
1588 Cypernsamtalen 1
1589 Cyprian 2
1590 D 2
1591 DA 12
1592 DB-datakälla 1
1593 DB-datakällor 1
1594 DDR 1
1595 DE 14
1596 DEBATT 2
1597 DISTINCT 1
1598 Da 3
1599 Dagen 1
1600 Dagens 8
1601 Dagerns 1
1602 Dagligen 3
1603 Dagmar 1
1604 Dagordningen 1
1605 Daily 1
1606 Dalai 7
1607 Dalmau 1
1608 Dam 3
1609 Damaskus 3
1610 Damer 1
1611 Dando 12
1612 Dandos 1
1613 Daniel 8
1614 Danmark 44
1615 Danmarks 2
1616 Danny 1
1617 Dansetteskivspelare 1
1618 Darmstadt 1
1619 Data 3
1620 Datablad 1
1621 Databladsläge 1
1622 Datum 1
1623 David 9
1624 Davids 1
1625 Davies 4
1626 Davis 2
1627 Dayton 2
1628 De 513
1629 Debatten 4
1630 Debatterna 1
1631 Decourrière 7
1632 Decourrièrebetänkandet 1
1633 Decourrières 3
1634 Definitionerna 1
1635 Definitivt 1
1636 Deklarationen 1
1637 Delat 1
1638 Delegationerna 1
1639 Dell'Alba 1
1640 Delningen 1
1641 Delors 8
1642 Delorskommissionens 1
1643 Delorsplanen 1
1644 Dels 2
1645 Deltagandet 1
1646 Delvis 2
1647 Dem 1
1648 Deminimus-bestämmelserna 1
1649 Demokrati 1
1650 Demokratiska 1
1651 Demonstranterna 1
1652 Den 626
1653 Denktash 2
1654 Denna 143
1655 Denne 1
1656 Deptford 1
1657 Deras 13
1658 Derbyshire 1
1659 Derivatmarknaden 1
1660 Derrick 1
1661 Desama 2
1662 Dess 7
1663 Dessa 123
1664 Dessutom 93
1665 Destabiliseringen 1
1666 Desto 3
1667 Det 2768
1668 Detaljerad 1
1669 Detaljerna 1
1670 Detaljområde 1
1671 Detektivbyrå 1
1672 Detsamma 3
1673 Detta 587
1674 Deutsche 3
1675 Devon 1
1676 Di 14
1677 Diagongränden 2
1678 Diagram 2
1679 Dialog 2
1680 Diamantopoulou 7
1681 Dig 1
1682 Digital 1
1683 Dimitrakopoulos 5
1684 Din 1
1685 Dineh 7
1686 Dinehbefolkningen 1
1687 Dinehindianerna 1
1688 Dior 1
1689 Dipecho 1
1690 Dipechos 2
1691 Diplomatiska 1
1692 Direktivet 18
1693 Direktivets 2
1694 Direktören 1
1695 Diskrimineringen 1
1696 Diskussionen 3
1697 Diskussionens 1
1698 Diskussionsämnet 1
1699 Diskuteras 1
1700 Dit 2
1701 Dixon 1
1702 Djupare 1
1703 Dobby 4
1704 Dobbys 1
1705 Dock 11
1706 Dokumenten 1
1707 Dokumentet 2
1708 Dom 4
1709 Domarna 1
1710 Dominique 3
1711 Domstolen 2
1712 Domstolens 2
1713 Don 9
1714 Donau 17
1715 Donaus 4
1716 Doris 2
1717 Dorothy 1
1718 Dos 3
1719 Doyles 1
1720 Doñana 2
1721 Doñana-katastrofen 1
1722 Dra 1
1723 Draco 8
1724 Drake 1
1725 Dricka 1
1726 Drive 5
1727 Drogheda 5
1728 Drug 1
1729 Dröjsmålet 1
1730 Du 47
1731 Dubbelt 1
1732 Dublin 5
1733 Dublinfonden 1
1734 Dublinkonventionen 2
1735 Dublinkonventionerna 1
1736 Dudley 19
1737 Dudleys 2
1738 Duhamels 1
1739 Duisenberg 3
1740 Duktig 1
1741 Dumbledore 1
1742 Dumpning 2
1743 Dunn 1
1744 Dupuis 4
1745 Dur 1
1746 Durban 1
1747 Dursley 9
1748 Dursleys 11
1749 Dutroux 1
1750 Dutroux-affären 1
1751 Dvs. 2
1752 Där 47
1753 Därav 4
1754 Därefter 13
1755 Däremot 26
1756 Därför 300
1757 Däri 1
1758 Därigenom 5
1759 Därmed 17
1760 Därtill 1
1761 Därute 1
1762 Därutöver 2
1763 Därvid 3
1764 Då 64
1765 Démocratique 1
1766 Díez 5
1767 Död 1
1768 Döda 2
1769 Dörrarna 1
1770 Dührkop 3
1771 E-kolibakteriesmittat 1
1772 ECB 2
1773 ECHO 13
1774 ECHO:s 1
1775 ECHR 2
1776 ECTAA 1
1777 EDD 3
1778 EDD-Gruppen 1
1779 EDD-gruppens 3
1780 EDF-medlens 1
1781 EDU:s 1
1782 EE 2
1783 EEC 1
1784 EEG 12
1785 EFTA:s 1
1786 EG 26
1787 EG-Israel 3
1788 EG-biståndet 1
1789 EG-direktiv 2
1790 EG-direktiven 2
1791 EG-direktivet 1
1792 EG-domstolen 25
1793 EG-domstolens 3
1794 EG-fördraget 9
1795 EG-kort 9
1796 EG-kortet 7
1797 EG-obligationer 1
1798 EG-rätt 2
1799 EG-rätten 1
1800 EG-verksamheter 1
1801 EG:s 8
1802 EIF 2
1803 EKSG 2
1804 EKSG-fördraget 6
1805 EL 9
1806 ELDR 3
1807 ELDR-gruppen 3
1808 ELDR:s 1
1809 EMU 3
1810 EMU-anpassningens 1
1811 EMU-anslutning 1
1812 EMU-eran 1
1813 EMU-fördraget 1
1814 EMU-kriterierna 2
1815 EMU-medlemsstater 1
1816 EMU-projekt 1
1817 EMU-projektet 1
1818 EMU-projektets 1
1819 EMU-samarbetet 1
1820 EMU:s 5
1821 EN 75
1822 ENS 10
1823 EPP-DE 1
1824 ERUF 1
1825 ES 7
1826 ETA 8
1827 ETA-förhandlare 1
1828 ETA:s 2
1829 EU 216
1830 EU- 2
1831 EU-AVS-avtalet 1
1832 EU-AVS-sammanhanget 1
1833 EU-Medelhavsområdet 1
1834 EU-anslutningen 1
1835 EU-behörighet 1
1836 EU-beslut 1
1837 EU-bistånd 1
1838 EU-biståndet 1
1839 EU-budgeten 1
1840 EU-enheten 1
1841 EU-fonder 1
1842 EU-fördrag 2
1843 EU-fördragen 1
1844 EU-fördraget 8
1845 EU-företag 2
1846 EU-förordningar 1
1847 EU-genomsnittet 1
1848 EU-initiativ 1
1849 EU-insatser 1
1850 EU-institutioner 1
1851 EU-institutionerna 4
1852 EU-institutionernas 2
1853 EU-kandidater 1
1854 EU-kommissionen 2
1855 EU-kort 2
1856 EU-kortet 2
1857 EU-kriterierna 1
1858 EU-lagstiftningen 4
1859 EU-landet 1
1860 EU-länder 7
1861 EU-länderna 6
1862 EU-ländernas 1
1863 EU-mantra 1
1864 EU-marknaden 1
1865 EU-marknader 1
1866 EU-medborgare 5
1867 EU-medborgarnas 1
1868 EU-medel 2
1869 EU-medlemmar 2
1870 EU-medlemmarna 2
1871 EU-medlemskap 2
1872 EU-medlemsstaterna 3
1873 EU-medlemsstaternas 1
1874 EU-miljöreglerna 1
1875 EU-nivå 6
1876 EU-nivån 1
1877 EU-ordförandeskapets 1
1878 EU-organ 2
1879 EU-pass 3
1880 EU-perspektiv 1
1881 EU-politik 1
1882 EU-program 2
1883 EU-regeringar 1
1884 EU-regi 1
1885 EU-reglerad 1
1886 EU-resurser 1
1887 EU-räntor 1
1888 EU-rätt 1
1889 EU-rättskipning 1
1890 EU-rådets 1
1891 EU-samarbetet 1
1892 EU-skeptiker 1
1893 EU-staterna 1
1894 EU-staternas 1
1895 EU-straffrätt 1
1896 EU-strukturfonder 1
1897 EU-system 1
1898 EU-sändebud 2
1899 EU-texterna 1
1900 EU-utvidgning 1
1901 EU-världen 1
1902 EU:s 125
1903 EUF 8
1904 EUF-medel 1
1905 EUF-medlen 1
1906 EUGFJ 4
1907 EUGFJ:s 1
1908 East 1
1909 Ecemis-förkastningslinjen 1
1910 Ecevit 2
1911 Echelon 3
1912 Echelon-nätet 1
1913 Edinburgh 3
1914 Editor 1
1915 Edward 1
1916 Edwards 3
1917 Effekten 3
1918 Effekterna 1
1919 Effektiv 2
1920 Effektiva 1
1921 Effektivitet 1
1922 Effektiviteten 2
1923 Eftarløn 2
1924 Efter 51
1925 Efterskalven 1
1926 Eftersom 73
1927 Efteråt 3
1928 Egeiska 1
1929 Egentligen 7
1930 Egypten 4
1931 Ehud 2
1932 Eichelberger 4
1933 Eichelbergers 1
1934 Eieck 1
1935 Ejido 26
1936 Ejidos 2
1937 Ekofin 2
1938 Ekofin-ministrar 1
1939 Ekofin-ministrarna 1
1940 Ekofin-rådet 8
1941 Ekologiskt 1
1942 Ekonomer 1
1943 Ekonomierna 1
1944 Ekonomin 4
1945 Ekonomisk 1
1946 Ekonomiska 6
1947 Ekonomistyrningen 1
1948 El 28
1949 Elbe 1
1950 Elden 1
1951 Elektriskt 1
1952 Elementen 1
1953 Elf 1
1954 Elfenbenskusten 1
1955 Elie 1
1956 Eline 1
1957 Elisabeth 1
1958 Eller 17
1959 Elles 3
1960 Elly 1
1961 Elmar 4
1962 Elorza 2
1963 Elst 1
1964 Elva 1
1965 Emellanåt 1
1966 Emellertid 12
1967 Emergency 1
1968 Emilia-Romagna 1
1969 Employment 1
1970 Employment-initiativen 1
1971 Emprego 1
1972 Empress 1
1973 En 282
1974 Enbart 1
1975 End 1
1976 Enda 1
1977 Endast 20
1978 Eneko 1
1979 Energisituationen 1
1980 Enfopol 1
1981 Engagemang 1
1982 Engelska 2
1983 Engelsmän 1
1984 England 10
1985 Englands 1
1986 Enigheten 1
1987 Enkelt 1
1988 Enligt 81
1989 Enorma 1
1990 Enrique 3
1991 Enterprise 1
1992 Entitet 1
1993 Equal 24
1994 Equal- 1
1995 Equal-betänkande 1
1996 Equal-betänkandet 10
1997 Equal-initiativet 19
1998 Equal-initiativets 2
1999 Equal-programmet 6
2000 Equal-programmets 1
2001 Equqal 2
2002 Er 8
2003 Era 4
2004 Erebus 1
2005 Erfarenheten 4
2006 Erfarenheter 1
2007 Erfarenheterna 4
2008 Ericsson 1
2009 Erika 44
2010 Erika-katastrofen 3
2011 Erika-katastrofer 1
2012 Erika-olyckan 1
2013 Erikas 14
2014 Erith 1
2015 Eritrea 1
2016 Erkki 2
2017 Ermua 1
2018 Eros 1
2019 Errols 1
2020 Ert 7
2021 Essen 1
2022 Essex 1
2023 Essex-Suffolk-Norfolkkusten 1
2024 Essexmaderna 1
2025 Estland 1
2026 Etiopien 5
2027 Etnisk 1
2028 Ett 149
2029 Etthundratjugotvå 1
2030 Euratom 4
2031 Euratomfördraget 1
2032 Euro 1
2033 Euro-Atlantiska 1
2034 Euro-Paper 1
2035 Euro-rådet 1
2036 Eurodac 4
2037 Eurodac-systemet 1
2038 Eurojust 6
2039 Euroland 3
2040 Euron 2
2041 Eurons 3
2042 Europa 710
2043 Europa-Afrika 1
2044 Europa-Medelhavsländerna 1
2045 Europademokrater 14
2046 Europademokraterna 2
2047 Europademokraternas 1
2048 Europadomstolen 1
2049 Europafrågan 1
2050 Europafrågor 1
2051 Europagrupp 1
2052 Europakonventionen 2
2053 Europaminister 2
2054 Europaministerns 1
2055 Europanivå 1
2056 Europaparlament 3
2057 Europaparlamentarikerna 1
2058 Europaparlamentet 288
2059 Europaparlamentets 118
2060 Europaparlamentsledamöternas 2
2061 Europarådet 2
2062 Europas 130
2063 Europaskatt 1
2064 Europatrupp 1
2065 Europaval 3
2066 Europavalen 4
2067 Europavalet 1
2068 Europavänligt 1
2069 Europe 4
2070 European 2
2071 Europeisk 1
2072 Europeiska 1197
2073 Europol 18
2074 Europolavtalet 1
2075 Europolkonventionen 1
2076 Europols 4
2077 Européerna 1
2078 Euroskeptikerna 1
2079 Eurostat 3
2080 Euskal 2
2081 Eusko 1
2082 Evans 7
2083 Evelyn 4
2084 Evelyns 1
2085 Eventuellt 2
2086 Exakt 1
2087 Excel 13
2088 Exceptionellt 1
2089 Exempel 6
2090 Exempelvis 2
2091 Exemplen 1
2092 Exemplet 2
2093 Experimental 1
2094 Experterna 3
2095 Expertutfrågningarna 1
2096 Explorer 2
2097 Exportera 6
2098 Expresso 1
2099 Extensible 3
2100 Exxon 3
2101 F 1
2102 F. 1
2103 FBI 2
2104 FEO 3
2105 FFP 1
2106 FFP:s 1
2107 FI 1
2108 FIPOL 1
2109 FMI 1
2110 FN 16
2111 FN-embargot 1
2112 FN-finansieringen 1
2113 FN-flyktingar 1
2114 FN-länder 1
2115 FN-närvaro 1
2116 FN-programmet 1
2117 FN-stadgan 1
2118 FN-stöd 1
2119 FN-uppdragets 1
2120 FN:s 36
2121 FPÖ 13
2122 FPÖ-ledaren 1
2123 FPÖ-medlemmar 1
2124 FPÖ:s 4
2125 FR 57
2126 FROM 1
2127 FRÅGOR 2
2128 FTSE 1
2129 FUF 1
2130 FYROM 8
2131 FYROM:s 4
2132 Fackföreningarna 1
2133 Fackföreningsrepresentanter 2
2134 Factortame-fallet 1
2135 Faim 1
2136 Fakta 2
2137 Faktum 12
2138 Fallet 5
2139 Falska 1
2140 Falskmyntning 1
2141 Falskt 1
2142 Falun 1
2143 Familjejordbruket 1
2144 Fan 1
2145 Far 9
2146 Farligt 1
2147 Farmor 5
2148 Farouk 1
2149 Fartyget 4
2150 Fartygets 1
2151 Fartygsbränslet 1
2152 Fascismen 1
2153 Faslane 2
2154 Faso 1
2155 Fast 7
2156 Fastän 1
2157 Fattas 1
2158 Fattigbasaren 1
2159 Fattigdomen 1
2160 Fattigdomsbekämpning 1
2161 Faulkner 2
2162 Federal 1
2163 Federation 1
2164 Feira 3
2165 Felaktigt 1
2166 Felet 1
2167 Fem 6
2168 Femte 1
2169 Femton 1
2170 Femårsprogrammet 1
2171 Ferber 1
2172 Fernando 5
2173 Fernández 4
2174 Ferte 1
2175 Festmåltider 1
2176 Festus 3
2177 Festus' 1
2178 Fidji-öarna 1
2179 Filen 1
2180 Filterfält 1
2181 Filtrera 4
2182 Filtrerad 1
2183 Filtrerat 1
2184 Filtreringsmetoder 1
2185 Fina 1
2186 Finansiella 1
2187 Finansiellt 1
2188 Finansiering 1
2189 Finansieringen 3
2190 Finansministrarna 1
2191 Finisterre 1
2192 Finland 27
2193 Finlands 1
2194 Finnarna 1
2195 Finner 2
2196 Finns 28
2197 Firman 1
2198 Fischler 18
2199 Fischlers 3
2200 Fishing 1
2201 Fisk 1
2202 Fiskare 1
2203 Fiskarnas 1
2204 Fiske 1
2205 Fiskeflottan 1
2206 Fiskeriförvaltning 3
2207 Fiskeriindustrin 1
2208 Fiskerisektorerna 1
2209 Fisket 2
2210 Fitousi 1
2211 Fitzsimons 1
2212 Fjolårets 1
2213 Fjorton 1
2214 Fjortonåriga 1
2215 Flandern 3
2216 Flautre 1
2217 Flautres 1
2218 Fleet 1
2219 Fleetwood 1
2220 Fler 2
2221 Flera 11
2222 Flertalet 1
2223 Flexibilitet 1
2224 Floden 2
2225 Floderna 1
2226 Flora 8
2227 Floras 1
2228 Florenz 19
2229 Florenzbetänkandet 1
2230 Flourish 1
2231 Flyg 1
2232 Flyg- 1
2233 Flygvärdinnorna 1
2234 Flytta 4
2235 Flyttfåglar 1
2236 Flämtande 1
2237 Flåsande 1
2238 Fléchard-affären 1
2239 FoU 1
2240 FoU-ramprogrammet 1
2241 Fodertillsatser 1
2242 Fog 1
2243 Folk 6
2244 Folkets 1
2245 Folkfronten 1
2246 Folkmordet 1
2247 Folkrepubliken 2
2248 Folkvalda 1
2249 Fondföretag 2
2250 Fondföretagen 1
2251 Fondsparande 1
2252 Fontaine 7
2253 Fontaines 1
2254 Food 1
2255 Force 1
2256 Ford 1
2257 Forestier 1
2258 Formulär 1
2259 Forskarna 1
2260 Forskningen 1
2261 Forsyth 1
2262 Forsyth-Byggen 1
2263 Fort 1
2264 Fortfarande 2
2265 Fortunas 1
2266 Fotografier 1
2267 Fraga 1
2268 Fraisse 1
2269 Fram 4
2270 Framför 11
2271 Framförallt 2
2272 Framgångarna 1
2273 Framläggandet 1
2274 Framsteg 1
2275 Framstegen 2
2276 Framställningar 1
2277 Framtagandet 1
2278 Framtida 1
2279 Framtiden 1
2280 Framåt 1
2281 France 2
2282 Frances 1
2283 Francis 3
2284 Franco 2
2285 Franklin 1
2286 Frankrike 63
2287 Frankrikes 10
2288 Franoise 1
2289 Fransmännen 3
2290 Franz 3
2291 François 1
2292 Frassoni 11
2293 Fred 19
2294 Freden 1
2295 Frederiksen 1
2296 Freds- 2
2297 Fredsprocessen 4
2298 Free 1
2299 Freetown 1
2300 Fricks 1
2301 Frid 1
2302 Frihet 3
2303 Friheten 1
2304 Frihetspartiet 3
2305 Frihetspartiets 1
2306 Fritt 1
2307 FrontPage 2
2308 Frontera 1
2309 Fru 213
2310 Fruteau 3
2311 Främjande 2
2312 Främjandet 1
2313 Främst 2
2314 Fråga 51
2315 Frågan 46
2316 Frågestund 4
2317 Frågor 6
2318 Frågorna 5
2319 Från 20
2320 Frånvaron 1
2321 Fukuyama 1
2322 Full 2
2323 Fund 4
2324 Fundera 1
2325 Fungerar 1
2326 Funktionen 1
2327 Fy 1
2328 Fyra 4
2329 Fyrtio 1
2330 Fysiska 1
2331 Fältpil 1
2332 Färden 1
2333 Färre 1
2334 Fästning 1
2335 Få 1
2336 Fågeln 1
2337 Får 16
2338 Följaktligen 8
2339 Följande 3
2340 Följden 3
2341 Följderna 2
2342 För 582
2343 Förbaskade 1
2344 Förbaskat 1
2345 Förbereda 1
2346 Förberedelserna 1
2347 Förbindelserna 1
2348 Förbrukningen 1
2349 Förbud 2
2350 Förbundskansler 1
2351 Förbundsrepubliken 5
2352 Fördelar 1
2353 Fördelarna 1
2354 Fördelen 2
2355 Fördomar 1
2356 Fördragen 2
2357 Fördraget 9
2358 Fördragets 1
2359 Före 8
2360 Förebyggande 2
2361 Föredragande 2
2362 Föredraganden 15
2363 Föredragandens 3
2364 Föredragningslista 3
2365 Föregående 1
2366 Förekommer 1
2367 Föreliggande 1
2368 Förenade 44
2369 Förenligheten 1
2370 Förenta 118
2371 Föresatsen 1
2372 Föreslagna 1
2373 Föreställer 1
2374 Föreställningen 1
2375 Företag 2
2376 Företrädaren 1
2377 Företrädarna 1
2378 Förfalskningar 1
2379 Förfarande 1
2380 Förfarandena 1
2381 Förfarandet 3
2382 Förflyttningen 1
2383 Förhandlingar 1
2384 Förhandlingen 1
2385 Förhindra 1
2386 Förhoppningar 1
2387 Förhoppningarna 2
2388 Förhoppningen 1
2389 Förhoppningsvis 4
2390 Förintelsekonferensen 1
2391 Förintelsen 2
2392 Förklaringen 1
2393 Förlisningen 1
2394 Förlorare 1
2395 Förlusterna 1
2396 Förlåt 2
2397 Förmodligen 3
2398 Förnyelsen 1
2399 Förordningen 4
2400 Förordningens 2
2401 Förorenaren 2
2402 Förpackningar 1
2403 Förr 1
2404 Förra 8
2405 Förresten 1
2406 Församlingarna 1
2407 Försiktighet 1
2408 Försiktighetsprincipen 2
2409 Förskjutningen 1
2410 Förslag 5
2411 Förslagen 5
2412 Förslaget 14
2413 Förslagets 1
2414 Förslagsrätt 1
2415 Först 60
2416 Första 3
2417 Förstainstansrätten 1
2418 Förstelning 1
2419 Förstå 1
2420 Förståeligt 1
2421 Förstår 3
2422 Förstörelsen 1
2423 Försvarsmakten 1
2424 Försämrar 1
2425 Försåvitt 1
2426 Försök 1
2427 Försöken 1
2428 Försöket 1
2429 Förtalet 1
2430 Förteckningen 2
2431 Förtjänster 1
2432 Förtroendet 1
2433 Förtrollad 1
2434 Förutom 13
2435 Förutsatt 2
2436 Förvaltningen 2
2437 Förvaltningsbolag 1
2438 Förvisso 5
2439 Förväntningarna 1
2440 Förvärrad 1
2441 Förändring 1
2442 Förändringar 3
2443 Förändringarna 2
2444 G8-mötet 1
2445 GA-stöd 1
2446 GAL 2
2447 GASP 1
2448 GATS-avtalen 1
2449 GATT 1
2450 GATT-avtalet 2
2451 GATT-förhandlingarna 1
2452 GATT:s 1
2453 GD 1
2454 GFP 1
2455 GJP 4
2456 GJP-reformerna 1
2457 GMO 16
2458 GMO-fri 1
2459 GRANT 1
2460 GUE 3
2461 GUSP 6
2462 GYLLENROY 1
2463 Gaeta 1
2464 Gai-Hinnom 4
2465 Galaprovinsen 1
2466 Galeote 4
2467 Galicien 6
2468 Gallagher 4
2469 Gallaghers 2
2470 Gallierna 1
2471 Gama 3
2472 Gamla 1
2473 Garanterandet 1
2474 García 1
2475 García-Margallo 2
2476 Garcías 1
2477 Gargani 5
2478 Gascognebukten 1
2479 Gasòliba 1
2480 Gatornas 1
2481 Gaulles 1
2482 Gaza 5
2483 Gazaregionen 1
2484 Gazaremsan 2
2485 Ge 1
2486 Gehenna 1
2487 Gemelli 1
2488 Gemensam 3
2489 Gemensamma 1
2490 Gemensamt 6
2491 Gemenskapen 1
2492 Gemenskapens 3
2493 Gemenskapsinitiativet 5
2494 Gemenskapsrätten 1
2495 Gemenskapsåtgärder 2
2496 Genast 1
2497 Gender 1
2498 Generaldirektorat 1
2499 Generaldirektoraten 1
2500 Generaldirektoratet 9
2501 Generaldirektören 1
2502 Generellt 1
2503 Genetiskt 2
2504 Genom 67
2505 Genomförande 1
2506 Genomförandet 4
2507 Genomsnittet 1
2508 Gentila 1
2509 Genua 1
2510 Genève 16
2511 Genèvekonventionen 7
2512 Genèvekonventionens 2
2513 Genèvekonventionerna 1
2514 Genèvemötet 1
2515 George 17
2516 Georgievski 1
2517 Ger 2
2518 Geremek 2
2519 Geresta 1
2520 Ghana 1
2521 Ghilardotti 1
2522 Gibraltar 1
2523 Gil-Delgado 1
2524 Gil-Robles 2
2525 Gillig 1
2526 Ginens 1
2527 Ginny 2
2528 Gino 1
2529 Giorgos 5
2530 Givet 1
2531 Givetvis 6
2532 Gjort 1
2533 Glansen 1
2534 Glase 1
2535 Glasgow 2
2536 Gligorov 1
2537 Global 1
2538 Globaliseringen 5
2539 Globaliseringens 1
2540 Glöm 1
2541 God 1
2542 Goddag 1
2543 Godkännandet 1
2544 Godspeed 1
2545 Goebbels 5
2546 Golan 6
2547 Golanhöjden 1
2548 Golanhöjderna 3
2549 Golden 1
2550 Golfströmmen 3
2551 Golgatavandring 1
2552 Gollnisch 2
2553 Gomes 1
2554 Gong-rörelsen 1
2555 González 2
2556 Goodwill 1
2557 Goodyear 14
2558 Gordon 1
2559 Gorka 1
2560 Gorostiaga 2
2561 Gorsel 3
2562 Gott 2
2563 Gouges 1
2564 Graal 1
2565 Graca 3
2566 Graco-affärerna 1
2567 Graefe 9
2568 Gran 1
2569 Granada 1
2570 Granger 5
2571 Grangers 1
2572 Granskningarna 1
2573 Granskningen 1
2574 Grants 1
2575 Grappakrigen 1
2576 Grattis 2
2577 Gratulerar 1
2578 Gravesend 1
2579 Gray's 1
2580 Graça 5
2581 Great 1
2582 Green 2
2583 Greenspan 1
2584 Greenwich 1
2585 Grekland 41
2586 Greklands 5
2587 Gringotts 4
2588 Grossetête 4
2589 Grosstête 1
2590 Grottor 1
2591 Group 1
2592 Grozny 3
2593 Grunden 4
2594 Grunderna 1
2595 Grundläggande 1
2596 Gruppen 42
2597 Grupperna 1
2598 Gruppnivåegenskaper 1
2599 Gryffindor 1
2600 Gränsarbetare 1
2601 Gränser 1
2602 Grått 1
2603 Gröna 3
2604 Gröner 2
2605 Grönitz 1
2606 Guatemala 1
2607 Gud 9
2608 Guds 3
2609 Guigou 1
2610 Guld- 1
2611 Guldsökare 1
2612 Gulfkriget 1
2613 Gulfområdet 1
2614 Gusp 1
2615 Guterres 11
2616 Guterrez 1
2617 Gutierres 1
2618 Gutíerrez 2
2619 Gwenzis 1
2620 Gyllenroy 3
2621 Gällande 1
2622 Gärna 1
2623 Gå 2
2624 Gång 2
2625 Går 1
2626 Gör 3
2627 Göra 1
2628 Göteborg 1
2629 Günther 1
2630 H-0002/99 1
2631 H-0006/00 1
2632 H-0020/00 1
2633 H-0021/00 1
2634 H-0022/00 1
2635 H-0024/00 1
2636 H-0025/00 1
2637 H-0026/00 1
2638 H-0027/00 1
2639 H-0028/00 1
2640 H-0029/00 1
2641 H-0031/00 1
2642 H-0035/00 1
2643 H-0036/00 1
2644 H-0040/00 1
2645 H-0041/00 1
2646 H-0042/00 1
2647 H-0044/00 1
2648 H-0045/00 1
2649 H-0045/99 1
2650 H-0049/00 1
2651 H-0052/00 1
2652 H-0053/00 1
2653 H-0057/00 1
2654 H-0095/00 1
2655 H-0117/00 1
2656 H-0122/00 1
2657 H-0209/99 1
2658 H-0218/97 1
2659 H-0237/97 1
2660 H-0778/99 1
2661 H-0780/99 1
2662 H-0781/99 1
2663 H-0782/99 1
2664 H-0785/99 1
2665 H-0786/99 1
2666 H-0788/99 1
2667 H-0791/99 1
2668 H-0793/99 1
2669 H-0795/99 1
2670 H-0796/99 1
2671 H-0798/99 1
2672 H-0801/99 1
2673 H-0805/99 1
2674 H-0807/99 1
2675 H-0808/99 1
2676 H-0813/99 1
2677 H-0817/99 1
2678 H-0819/99 1
2679 H-0829/99 1
2680 H. 1
2681 H.C. 1
2682 HELP 1
2683 HON 1
2684 HOTREC 1
2685 HTML 2
2686 HTML-formatet 1
2687 HTML-kod 1
2688 Haag 3
2689 Haarder 5
2690 Habana 1
2691 Habitat 1
2692 Hade 4
2693 Hadera 1
2694 Hagrid 7
2695 Hague 1
2696 Haider 26
2697 Haiderpolitiken 1
2698 Haiders 24
2699 Haifa 1
2700 Hain 1
2701 Hainaut 1
2702 Halonen 1
2703 Halva 1
2704 Hamburg 2
2705 Hamilton 1
2706 Hamna 1
2707 Hamnarna 1
2708 Hamnens 1
2709 Han 295
2710 Handeln 1
2711 Handelsavtal 1
2712 Handelsavtalet 1
2713 Handikappades 1
2714 Handikapporganisationer 1
2715 Handlingen 1
2716 Handlingskraften 1
2717 Hangarfartyget 1
2718 Hans 19
2719 Hanteringen 1
2720 Har 31
2721 Harbour 2
2722 Harbours 1
2723 Harmoniseringsbyrån 1
2724 Harold 1
2725 Harry 116
2726 Harrys 14
2727 Harwich 1
2728 Hatzidakis 3
2729 Hatzidakisbetänkandet 1
2730 Haug 1
2731 Hautala 4
2732 Havel 10
2733 Havels 2
2734 Haven 1
2735 Havet 1
2736 Havsprodukternas 1
2737 Havsvärlden 1
2738 Heathrow 2
2739 Heaton-Harris 1
2740 Hebreiska 1
2741 Hebriderna 1
2742 Hebron- 1
2743 Hecke 3
2744 Heckes 2
2745 Hedge 1
2746 Hedkvist 1
2747 Hedwig 5
2748 Hedwigs 2
2749 Hefaistos 1
2750 Heidi 1
2751 Heights 1
2752 Heinz 1
2753 Hej 2
2754 Hela 14
2755 Helighet 1
2756 Helmkom-avtalet 1
2757 Helms-Burton 1
2758 Help 1
2759 Helsingfors 52
2760 Helsingfors-besluten 1
2761 Helsingforskonventionen 1
2762 Helsingforsmandatet 1
2763 Helsingforsmötet 2
2764 Helsingforstoppmötet 1
2765 Helt 8
2766 Hemliga 1
2767 Hemma 1
2768 Hennes 9
2769 Henry 2
2770 Herman 1
2771 Hermes 1
2772 Hermione 10
2773 Hernandez 1
2774 Hernández 1
2775 Herr 965
2776 Herre 1
2777 Herregud 1
2778 Herritarrok 2
2779 Hertfordshire 1
2780 Hicks 1
2781 Hilton 1
2782 Himalaya 1
2783 Himalayabergen 1
2784 Hind 1
2785 Hinken 1
2786 Hinner 1
2787 Historien 6
2788 Hit 4
2789 Hitler 8
2790 Hitler-regimen 1
2791 Hitlers 1
2792 Hittills 8
2793 Hjalmar 8
2794 Hjälp 3
2795 Hoechst 1
2796 Hogwarts 12
2797 Holland 3
2798 Hollywoodfilmer 1
2799 Holzmann 1
2800 Holzmann-gruppen 1
2801 Hon 75
2802 Honduras 2
2803 Hong 1
2804 Hongkong 4
2805 Hoogoven 1
2806 Hoppet 2
2807 Horizon 2
2808 Horst 1
2809 Hos 1
2810 Hotel 5
2811 Hotelsemönstret 1
2812 Hoti 1
2813 House 1
2814 Howard 1
2815 Howittsbetänkandet 1
2816 Hubert 1
2817 Hudghton 8
2818 Hudghtons 1
2819 Hudsonfloden 1
2820 Hugg 1
2821 Hughes 1
2822 Huhne 5
2823 Huj 4
2824 Hulten 12
2825 Hultenbetänkandet 4
2826 Hultens 3
2827 Hulthen 4
2828 Hulthens 2
2829 Human 1
2830 Hun 1
2831 Hundratals 1
2832 Hungersnöd 1
2833 Hur 116
2834 Hurdana 1
2835 Huruvida 3
2836 Huset 1
2837 Hustrun 2
2838 Huvudaktörerna 1
2839 Huvudansvaret 1
2840 Huvudbudskapet 1
2841 Huvuddelen 1
2842 Huvudfrågorna 1
2843 Huvudlinjen 1
2844 Huvudmålet 1
2845 Huvudmålsättningen 1
2846 Huvudproblemet 1
2847 Huvudregeln 1
2848 Huvudsaken 3
2849 Hyckleri 1
2850 Häkkinens 1
2851 Häktningsorder 1
2852 Hälften 1
2853 Händelsen 1
2854 Händelser 1
2855 Händelserna 3
2856 Hängde 1
2857 Hänsch 2
2858 Hänsyn 3
2859 Här 86
2860 Härav 2
2861 Härigenom 1
2862 Härmed 6
2863 Härom 1
2864 Häromdagen 1
2865 Hästen 2
2866 Håll 3
2867 Hållbar 2
2868 Håller 1
2869 Hög 3
2870 Höga 1
2871 Höge 1
2872 Högerextremism 1
2873 Högnivågruppen 2
2874 Högre 1
2875 Högst 1
2876 Högvärdighet 1
2877 Höjden 1
2878 Hör 1
2879 I 888
2880 I-programmet 2
2881 I. 1
2882 IBM 1
2883 ICCAT 6
2884 ICCAT:s 2
2885 ICES 1
2886 ICES-zon 1
2887 ICES-zonen 1
2888 ICES-zonerna 1
2889 ICT-företag 1
2890 IDEA-åldern 1
2891 IFOP 1
2892 IGC 4
2893 II 28
2894 II-programmet 4
2895 III 26
2896 III- 1
2897 III-gränser 1
2898 III-initiativet 1
2899 III-programmet 2
2900 IIIA 1
2901 IIIC 2
2902 ILA 21
2903 ILO 2
2904 IMF 1
2905 IMO 2
2906 IMO:s 1
2907 INTE 1
2908 INTERREG 2
2909 INTERREG-initiativ 1
2910 IOPCF 2
2911 IOPCF:s 1
2912 IRA 1
2913 ISA 1
2914 ISD 1
2915 ISPA-instrumentet 1
2916 IT 9
2917 IT-branschen 1
2918 IT-fattiga 1
2919 IT-infrastruktur 2
2920 IT-rika 1
2921 IT-utvecklingen 1
2922 ITALIENSKA 1
2923 IV 5
2924 IX 2
2925 Ibland 8
2926 Icke 5
2927 Icke-statliga 1
2928 Idén 3
2929 Igal 1
2930 Igår 1
2931 Ihållande 1
2932 Ikväll 1
2933 Ile-de-France 1
2934 Ilisu- 1
2935 Ilisudammen 4
2936 Illa 1
2937 Illegalt 1
2938 Ilsket 1
2939 Imbeni 3
2940 Immigrationen 1
2941 Importera 1
2942 Inbillar 1
2943 Inbördes 1
2944 Indien 6
2945 Indiens 1
2946 Indikatorerna 1
2947 Indirekt 1
2948 Indiska 1
2949 Indonesien 11
2950 Industriella 1
2951 Industrin 1
2952 Industrins 1
2953 Infektiös 1
2954 Information 2
2955 Informationen 2
2956 Informationscentren 1
2957 Informationssamhället 1
2958 Infödingsmattor 1
2959 Inför 10
2960 Införandet 4
2961 Inga 8
2962 Ingen 29
2963 Ingenstans 2
2964 Ingenting 5
2965 Inger 1
2966 Inget 9
2967 Ingetdera 1
2968 Inglewood 1
2969 Inglewoods 1
2970 Ingusjien 1
2971 Initiativ 1
2972 Initiativet 6
2973 Initiativets 1
2974 Inklusive 1
2975 Inkomstklyftan 1
2976 Inlåst 1
2977 Inlåsta 1
2978 Inn 1
2979 Innan 20
2980 Innebär 1
2981 Innebörden 1
2982 Innehållet 1
2983 Innehållsmässigt 1
2984 Innovation 1
2985 Inom 30
2986 Inre 2
2987 Inresan 1
2988 Inriktning 1
2989 Inrättandet 1
2990 Insamling 1
2991 Insatserna 2
2992 Insatsstyrkan 1
2993 Inskränkningarna 1
2994 Insolvens 1
2995 Insolvensförfaranden 1
2996 Installera 1
2997 Institute 1
2998 Institutionellt 1
2999 Instrumenten 2
3000 Inte 63
3001 Integra 2
3002 Integritet 1
3003 Intellectual 2
3004 Intern 1
3005 International 7
3006 Internationell 2
3007 Internationella 24
3008 Internet 40
3009 Internet-ekonomins 1
3010 Internetrevolutionen 2
3011 Internetrevolutionens 1
3012 Interreg 71
3013 Interreg- 1
3014 Interreg-anslag 1
3015 Interreg-anslagen 1
3016 Interreg-initiativ 1
3017 Interreg-initiativet 9
3018 Interreg-programmen 1
3019 Interreg-programmet 2
3020 Interreg-riktlinjer 1
3021 Interreg-ärendena 1
3022 Interregs 4
3023 Interventionspriser 1
3024 Intill 2
3025 Intressant 1
3026 Invandrarna 1
3027 Investeringar 2
3028 Investeringsnivåerna 1
3029 Investments 1
3030 Irak 5
3031 Iraks 1
3032 Iran 3
3033 Irans 1
3034 Irland 52
3035 Irlands 2
3036 Irländska 7
3037 Isabel 3
3038 Island 1
3039 Isler 2
3040 Ismail 1
3041 Isoza-floden 1
3042 Ispa 1
3043 Ispa- 1
3044 Ispar 1
3045 Israel 81
3046 Israel-Syrienfrågan 1
3047 Israeliska 1
3048 Israelkritik 1
3049 Israels 18
3050 Istanbul 1
3051 Istället 3
3052 Italien 40
3053 Italiens 1
3054 Ivanov 1
3055 Izquierdo 1
3056 J 3
3057 JAG 1
3058 Ja 55
3059 Ja-så-är-vi-här-igen-leende 1
3060 Jackson 2
3061 Jacob 2
3062 Jacques 8
3063 Jaffa 2
3064 Jag 2866
3065 Jaga 1
3066 Jaha 2
3067 Jakov 1
3068 Jamaica 2
3069 Jamen 3
3070 James 5
3071 Jan 3
3072 Jan-Kees 1
3073 Japan 9
3074 Jarzembowski 3
3075 Jaså 5
3076 Javette-Le 1
3077 Javier 9
3078 Jean 5
3079 Jean-Claude 2
3080 Jean-Olivier 1
3081 Jefferson 1
3082 Jens-Peter 1
3083 Jeremia 1
3084 Jersey 2
3085 Jerusalem 12
3086 Jerusalems 4
3087 Jesus 1
3088 Jet 1
3089 Jo 8
3090 Jo-Ann 2
3091 Joakim 1
3092 Joaquim 1
3093 Joaquín 1
3094 Jobs 2
3095 Jodå 1
3096 Johan 1
3097 John 17
3098 Jojon 2
3099 Jomän 1
3100 Jonas 2
3101 Jonckheer 9
3102 Jonckheerbetänkandet 3
3103 Jonckheers 3
3104 Jord 1
3105 Jordan 1
3106 Jordanien 1
3107 Jordanierna 1
3108 Jordans 1
3109 Jordbruk 2
3110 Jordbrukande 1
3111 Jordbruket 3
3112 Jordbruksekonomin 1
3113 Jordbruksministeriet 1
3114 Jorge 3
3115 Josafats 1
3116 Joseph 1
3117 Jospin 3
3118 José 2
3119 Journal 1
3120 Journalisten 1
3121 Journalister 2
3122 Journalists 1
3123 Jove 4
3124 Jovisst 1
3125 Joyces 1
3126 Ju 6
3127 Judarna 1
3128 Judegrabbens 1
3129 Jugoslavien 32
3130 Jugoslaviens 7
3131 Juncker 1
3132 Junker 1
3133 Junkers 1
3134 Juridisk 1
3135 Just 35
3136 Justering 7
3137 Justeringen 1
3138 Jämförelse 1
3139 Jämfört 4
3140 Jämställdhet 2
3141 Jämställdheten 1
3142 Jämställdhetsaspekter 1
3143 Jörg 18
3144 Jösses 2
3145 Júcar 2
3146 KFOR 1
3147 KLM 1
3148 KOM(1997 1
3149 KOM(1998 5
3150 KOM(1999 21
3151 KOM(1999)0003 2
3152 KOM(1999)0598 1
3153 KOM(98)0662 1
3154 KOM(99)0598 1
3155 Kabila 1
3156 Kabul 1
3157 Kackerlackor 1
3158 Kafferast 1
3159 Kafor 1
3160 Kairo 2
3161 Kaleidoskop 2
3162 Kalejdoskop 1
3163 Kambodja 14
3164 Kambodjas 1
3165 Kammaren 5
3166 Kampen 1
3167 Kan 53
3168 Kanada 6
3169 Kanarieöarna 2
3170 Kandalprovinsen 1
3171 Kandidatländerna 1
3172 Kandidatländernas 1
3173 Kano 1
3174 Kanske 20
3175 Kantabrien 3
3176 Kapital- 1
3177 Kaptenen 1
3178 Karamanous 1
3179 Karas 4
3180 Karelen 1
3181 Karibien 5
3182 Karin 1
3183 Karl 6
3184 Karl-Heinz 2
3185 Karlsruhe 2
3186 Kartellamt 1
3187 Kartellförbudet 1
3188 Kaspiska 1
3189 Katalonien 1
3190 Katastrofen 1
3191 Katastrofer 1
3192 Kategorifältområde 1
3193 Katiforis 26
3194 Katiforisbetänkandet 2
3195 Kaufmann 1
3196 Kaukasus 4
3197 Kauppi 2
3198 Kazakstan 1
3199 Kedourie 3
3200 Kedouries 1
3201 Kejsarens 1
3202 Kennedy 1
3203 Kensington 1
3204 Kente 2
3205 Kenyatta 1
3206 Kermit 1
3207 Kfor 1
3208 Kfor-styrkan 1
3209 Kfor-styrkorna 1
3210 Kfor-trupperna 1
3211 Khartum 1
3212 Khatami 2
3213 Kina 44
3214 Kinapolitik 1
3215 Kinas 4
3216 Kindermann 3
3217 Kinnock 29
3218 Kinnocks 5
3219 Kirgizistan 5
3220 Kit 1
3221 Kjolarna 1
3222 Klart 1
3223 Klimas 1
3224 Klippan 1
3225 Klistra 1
3226 Klockan 4
3227 Knappt 1
3228 Knörr 7
3229 Koch 15
3230 Kochs 1
3231 Kocken 1
3232 Kod 1
3233 Koden 1
3234 Kofi 1
3235 Kohl 1
3236 Kohoutek 1
3237 Kollega 1
3238 Kollegan 3
3239 Kolleger 3
3240 Kollektiva 1
3241 Kom 7
3242 Kommer 33
3243 Kommissarie 1
3244 Kommissionen 202
3245 Kommissionens 62
3246 Kommissionsledamöterna 1
3247 Kommissionär 22
3248 Kommissionären 9
3249 Kommissionärerna 1
3250 Kommittologi 1
3251 Kommittéförfarande 2
3252 Kommitténs 1
3253 Kommuner 1
3254 Kommunerna 1
3255 Kompletterande 1
3256 Kompromissformuleringar 1
3257 Koncentrationen 1
3258 Konceptet 2
3259 Konflikten 2
3260 Kongo 6
3261 Kongressen 1
3262 Kongs 1
3263 Konkret 1
3264 Konkreta 1
3265 Konkurrens 3
3266 Konkurrensen 6
3267 Konkurrenspolitik 1
3268 Konkurrenspolitiken 4
3269 Konkurrensprincipen 2
3270 Konrad 1
3271 Konsekvenserna 3
3272 Konstigt 1
3273 Konsumenten 1
3274 Konsumenterna 4
3275 Konsumentpolitiken 1
3276 Kontoren 1
3277 Kontroll 1
3278 Kontroller 4
3279 Kontrollfunktionen 1
3280 Kontrollförfarandet 1
3281 Kontrollnamn 1
3282 Kontrollstöd 1
3283 Konventionen 4
3284 Konventioner 1
3285 Konvertera 1
3286 Kopiera 3
3287 Kopplat 1
3288 Korea 3
3289 Korrekt 1
3290 Korridorerna 1
3291 Kors 1
3292 Korsfrågor 1
3293 Kort 11
3294 Kortfattat 2
3295 Koschermat 1
3296 Kososvokonflikten 1
3297 Kosova 1
3298 Kosovo 176
3299 Kosovoalbanerna 1
3300 Kosovofrågan 1
3301 Kosovoinsatser 1
3302 Kosovokonflikten 3
3303 Kosovokriget 2
3304 Kosovokrigets 1
3305 Kosovoproblemet 1
3306 Kosovos 17
3307 Kostnaden 1
3308 Kostnaderna 5
3309 Kotka 1
3310 Kouchener 1
3311 Kouchner 14
3312 Kouchners 9
3313 Koushner 1
3314 Koushners 2
3315 Kraftiga 1
3316 Krajina 1
3317 Krav 1
3318 Kraven 1
3319 Kravet 2
3320 Kreml 1
3321 Kriget 3
3322 Krigsherrar 1
3323 Kriterier 1
3324 Kroatien 6
3325 Kronos 1
3326 Kroppen 1
3327 Kuba 22
3328 Kubas 6
3329 Kuckelkorn 1
3330 Kultur 20
3331 Kulturell 3
3332 Kulturellt 1
3333 Kulturen 1
3334 Kumar 1
3335 Kunde 1
3336 Kunder 2
3337 Kundorder 1
3338 Kungliga 1
3339 Kunskapssamhället 1
3340 Kurti 1
3341 Kurtz 7
3342 Kusligt 1
3343 Kuwait 1
3344 Kv3 1
3345 Kvalitet 2
3346 Kvalitén 1
3347 Kvantifierade 1
3348 Kvartal 1
3349 Kvestorerna 1
3350 Kvicksilver 1
3351 Kvinnan 2
3352 Kvinnor 22
3353 Kvinnorna 7
3354 Kvinnornas 4
3355 Kvinnors 2
3356 Kvotering 1
3357 Kväkareuropa 1
3358 Kyi 1
3359 Kyoto 6
3360 Kyoto-protokollet 1
3361 Kyotoprocesserna 1
3362 Kyotoprotokollet 2
3363 Kyotos 1
3364 Kypare 1
3365 Känner 4
3366 Känsliga 1
3367 Kära 16
3368 Käraste 1
3369 Käre 1
3370 Kärnan 1
3371 Kärnkraftverk 1
3372 Kärnkraftverket 1
3373 Kärnten 3
3374 Köhler 1
3375 Köket 1
3376 Köln 7
3377 Kölnprocessen 2
3378 Kön 1
3379 Köpenhamn 4
3380 L 1
3381 LEVE 1
3382 LIMIT 1
3383 LOCKMAN 1
3384 LTCM 1
3385 La 8
3386 Laan 2
3387 Laans 5
3388 Labourregeringens 1
3389 Labours 1
3390 Lagkatalogen 1
3391 Lagstiftningen 1
3392 Lama 5
3393 Lamas 2
3394 Lancker 3
3395 Land 1
3396 Landaburu 1
3397 Landet 4
3398 Landis 1
3399 Landsbygden 1
3400 Landsbygdens 1
3401 Landsbygdsområdena 1
3402 Lange 12
3403 Langen 13
3404 Langenbetänkandet 1
3405 Langens 3
3406 Langer 2
3407 Langes 1
3408 Language 3
3409 Lanka 3
3410 Lannoye 4
3411 Lannoyes 1
3412 Lappland 3
3413 Lapus 1
3414 Larcher 1
3415 Lastbilen 1
3416 Lastbilstrafiken 1
3417 Lasten 1
3418 Latina 2
3419 Latinamerika 1
3420 Laurent 1
3421 Le 4
3422 Leader 47
3423 Leader+ 25
3424 Leader+-initiativen 1
3425 Leader+-programmen 1
3426 Leader+-programmet 6
3427 Leader-initiativet 3
3428 Leader-programmen 1
3429 Leader-programmens 1
3430 Leader-programmet 4
3431 Leader-projekten 1
3432 Leader-stödområdena 1
3433 Lechner 2
3434 Leclerc 1
3435 Ledamot 4
3436 Ledamoten 7
3437 Ledamotens 1
3438 Ledamöter 4
3439 Ledamöterna 2
3440 Ledare 1
3441 Ledningen 1
3442 Lee 1
3443 Leendet 1
3444 Legenden 2
3445 Leinemanns 2
3446 Leinen 7
3447 Leinens 1
3448 Leinster 1
3449 Leinsters 1
3450 Leonardo 1
3451 Leone 1
3452 Leoni 1
3453 Lepos 1
3454 Lesotho 1
3455 Lettland 1
3456 Levande 1
3457 Levante 1
3458 Libanon 6
3459 Liberal 2
3460 Liberaliseringen 1
3461 Liberty 2
3462 Libyens 1
3463 License 1
3464 Lider 1
3465 Lieneman 1
3466 Lienemann 19
3467 Lienemannbetänkandet 1
3468 Lienemanns 9
3469 Lienemannsbetänkandet 1
3470 Life 52
3471 Life-Miljö 1
3472 Life-Natur 1
3473 Life-Tredje 1
3474 Life-förordningen 1
3475 Life-instrumentet 1
3476 Life-miljö 1
3477 Life-natur 1
3478 Life-programmen 1
3479 Life-programmet 2
3480 Life-programmets 1
3481 Life-projekt 1
3482 Life-projektets 1
3483 Life:s 2
3484 Lifes 1
3485 Liikanen 14
3486 Lika 1
3487 Likadant 1
3488 Likafullt 2
3489 Likaså 6
3490 Like 1
3491 Liknande 1
3492 Likriktning 1
3493 Liksom 17
3494 Likväl 4
3495 Lille 1
3496 Lillehammer-rapporten 1
3497 Limpopodalen 1
3498 Lindgren 2
3499 Linds 1
3500 Link 1
3501 Links 1
3502 Lipietz 1
3503 Lissabon 83
3504 Lissabon-initiativ 1
3505 Lissabonmötet 4
3506 Listorna 1
3507 Litauen 3
3508 Lite 1
3509 Litteraturen 1
3510 Little 1
3511 Liverpool 3
3512 Livliga 9
3513 Livsmedelssäkerhet 2
3514 Livsmedelssäkerheten 2
3515 Livsmedelssäkerhetsmyndigheten 1
3516 Livsmedelssäkerhetsprogram 1
3517 Livsmedelsäkerhet 1
3518 Ljuden 1
3519 Ljug 1
3520 Ljuspunkterna 1
3521 Lloyds 1
3522 Lockman 3
3523 Lockmans 1
3524 Logiskt 1
3525 Loi 1
3526 Loire 1
3527 Loire-Atlantique 2
3528 Lokala 1
3529 Lomas 1
3530 Lomé 3
3531 Loméavtal 1
3532 Loméavtalens 1
3533 Loméavtalet 2
3534 Lomékonvention 1
3535 Lomékonventionen 18
3536 Lomékonventionens 3
3537 Lomékonventionerna 1
3538 Loméländerna 1
3539 Lomémodellen 1
3540 Loméramen 1
3541 Lomésamarbetet 1
3542 Loméuppgörelse 1
3543 London 15
3544 Lord 4
3545 Lorenzettis 1
3546 Lorosae 1
3547 Lorraine 2
3548 Lothar 3
3549 Louis 4
3550 Lousewies 1
3551 Louth 1
3552 Loyola 2
3553 Lucas 6
3554 Lucius 1
3555 Luften 2
3556 Lugard 1
3557 Luis 2
3558 Lukten 1
3559 Lulling 2
3560 Luncheonette 1
3561 Lund 2
3562 Luren 1
3563 Lutte 1
3564 Luxemburg 21
3565 Luxemburgprocess 3
3566 Luxemburgprocessen 6
3567 Luxemburgprocessens 1
3568 Luxemburgs 1
3569 Luxemburgstrategin 1
3570 Lycka 1
3571 Lyckas 1
3572 Lyckligt- 1
3573 Lyckligtvis 4
3574 Lyncharna 1
3575 Lynne 2
3576 Lynnes 2
3577 Lyon 1
3578 Lyssna 1
3579 Läget 3
3580 Lägg 7
3581 Lägga 2
3582 Lägre 1
3583 Lämna 1
3584 Lämplig 1
3585 Lämpliga 1
3586 Lämpligt 1
3587 Länder 2
3588 Längs 1
3589 Länka 2
3590 Lärande 1
3591 Läs 3
3592 Lån 1
3593 Långrandigt 1
3594 Långsamheten 1
3595 Långt 1
3596 Låt 149
3597 Lönsamhet 1
3598 Lösningarna 1
3599 Lösningen 3
3600 Lööw 2
3601 Lübeck 1
3602 MARPOL 1
3603 MATEN 1
3604 MPLA 2
3605 MSDN 1
3606 MSF 1
3607 Maaaaaammma 1
3608 Maastricht 4
3609 Maastrichtfördraget 7
3610 Maastrichtkonferensen 1
3611 Maastrichtkriterierna 2
3612 Maaten 3
3613 MacCormick 6
3614 Macao 2
3615 Mace 1
3616 Machie 1
3617 Madagaskar 2
3618 Madeira 3
3619 Madison 2
3620 Madrid 4
3621 Madrid- 1
3622 Maes 6
3623 Maghreb 1
3624 Maghrebländerna 1
3625 Maij-Weggen 4
3626 Maij-Weggens 1
3627 Mainstreaming 1
3628 Majestäts 1
3629 Major 1
3630 Majoriteten 3
3631 Makedonien 66
3632 Makedoniens 5
3633 Makten 1
3634 Maktproblem 1
3635 Malfoy 14
3636 Malfoys 1
3637 Mallorca 1
3638 Malmström 3
3639 Malone 1
3640 Malta 42
3641 Maltas 4
3642 Mamma 1
3643 Mamère 1
3644 Man 195
3645 Managing 1
3646 Manchester 2
3647 Mandela 1
3648 Mandelstam 2
3649 Manhattan 1
3650 Mannen 5
3651 Manuel 1
3652 Manyema 1
3653 Mappen 1
3654 Maputo 1
3655 Marches 1
3656 Mare 1
3657 Margarin 1
3658 Marginaliseringen 1
3659 Margot 11
3660 Maria 2
3661 Marie 1
3662 Marie-Noëlle 2
3663 Marindepartementet 1
3664 Marinho 5
3665 Marinhos 1
3666 Mario 2
3667 Maritain 1
3668 Markera 1
3669 Marknaden 4
3670 Marknadsverkan 1
3671 Markov 4
3672 Marlow 4
3673 Marlows 1
3674 Marocko 7
3675 Marpol-fördraget 1
3676 Marpolkonventionen 2
3677 Marques 1
3678 Marseille 1
3679 Marset 1
3680 Marshallplan 1
3681 Marshallplanen 1
3682 Marshallplaner 1
3683 Martin 4
3684 Martinez 2
3685 Martini 1
3686 Martín 4
3687 Martíns 1
3688 Masker 1
3689 Mason 3
3690 Massor 1
3691 Matematiker 1
3692 Mathieu 1
3693 Matisse 1
3694 Matrovica 1
3695 Matrovicas 1
3696 Max 1
3697 Maximalt 1
3698 Maximiåldern 1
3699 McCarthy 7
3700 McCartin 1
3701 McGowan 1
3702 McKenna 2
3703 McNally 3
3704 McNallybetänkandet 1
3705 McNallys 1
3706 Meat 1
3707 Mebeki 1
3708 Med 148
3709 Meda 7
3710 Meda-programmet 2
3711 Medan 27
3712 Medbeslutande 1
3713 Medborgare 2
3714 Medborgaren 1
3715 Medborgarna 7
3716 Medborgarnas 1
3717 Meddelande 1
3718 Medel 1
3719 Medelhavet 22
3720 Medelhavets 5
3721 Medelhavshamnar 2
3722 Medelhavsländer 1
3723 Medelhavsländerna 5
3724 Medelhavsområdet 8
3725 Medelhavsområdets 1
3726 Medelhavsregionen 2
3727 Medelhavstonfisken 1
3728 Medellängd 1
3729 Medger 1
3730 Medicinen 1
3731 Medina 5
3732 Medlemsstaterna 12
3733 Medlemsstaternas 3
3734 Medresenärerna 1
3735 Medvetandet 1
3736 Meijer 1
3737 Mekanisk 1
3738 Mellan 5
3739 Mellanöstern 44
3740 Mellanösternfreden 1
3741 Mellanösterns 2
3742 Memoirs 1
3743 Men 601
3744 Menar 2
3745 Meningen 2
3746 Mentaliteten 1
3747 Menéndez 1
3748 Mer 19
3749 Merseybeat 1
3750 Messias 1
3751 Mest 1
3752 Metallräcket 1
3753 Metis 3
3754 Mets 4
3755 Mexico 1
3756 Mexiko 3
3757 Michel 5
3758 Michelin 4
3759 Michelin-koncernen 1
3760 Michiel 1
3761 Microsoft 29
3762 Middelhoek 1
3763 Midlands 2
3764 Miert 1
3765 Mika 1
3766 Milano 1
3767 Milano-området 1
3768 Miles 1
3769 Militär 1
3770 Miljoner 1
3771 Miljöaspekterna 1
3772 Miljöinstitutioner 1
3773 Miljökatastrof 1
3774 Miljökatastrofen 1
3775 Miljökatastroferna 1
3776 Miljömässigt 1
3777 Miljön 2
3778 Miljöproblem 1
3779 Miljöproblemen 1
3780 Miljösituationen 1
3781 Miljövariabeln 1
3782 Millennierundan 1
3783 Millennium 3
3784 Miller 3
3785 Milosevic 11
3786 Milosevic-regimen 1
3787 Milosevicregimen 1
3788 Milosevics 6
3789 Min 114
3790 Mina 35
3791 Minchah-bön 1
3792 Mindre 2
3793 Minimiregler 1
3794 Minimistorleken 1
3795 Minister 1
3796 Ministeriet 3
3797 Ministern 2
3798 Ministerrådet 1
3799 Minnen 1
3800 Minnesota 1
3801 Minns 2
3802 Minoriteter 1
3803 Minsk 1
3804 Minskar 1
3805 Minskningen 1
3806 Minst 1
3807 Minsta 1
3808 Minuc 1
3809 Mira 2
3810 Mirakel 1
3811 Miranda 1
3812 Mishkenot 1
3813 Mississippi 2
3814 Mister 2
3815 Mitrovic 1
3816 Mitrovica 17
3817 Mitt 20
3818 Mitterrand 1
3819 Mitterrands 1
3820 Moabs 1
3821 Mobiliseringen 1
3822 Moder 2
3823 Modern 1
3824 Modernare 1
3825 Modernisering 1
3826 Modrow 1
3827 Mohieddin 1
3828 Moldavien 1
3829 Mollar 2
3830 Molly 3
3831 Moloksdyrkarna 1
3832 Moluckerna 3
3833 Mom's 1
3834 Monde 3
3835 Mongoliet 2
3836 Monica 1
3837 Monika 2
3838 Monnet 1
3839 Monnets 1
3840 Monsieur 1
3841 Montego 1
3842 Montenegro 2
3843 Monti 28
3844 Monti-paketet 1
3845 Montipaketet 1
3846 Montis 1
3847 Montreal 4
3848 Mor 7
3849 Moral 1
3850 Moratinos 4
3851 Moratorium 1
3852 Morbihan 1
3853 Morbror 5
3854 Morgan 6
3855 Morgantini 5
3856 Morgantinis 1
3857 Morillon 2
3858 Morse 1
3859 Moseboken 1
3860 Moses 1
3861 Moshe 1
3862 Moskva 3
3863 Moss 1
3864 Moster 2
3865 Mot 25
3866 Motiveringen 1
3867 Motorn 1
3868 Motsättningar 1
3869 Mottagningsanordningar 1
3870 Mount 1
3871 Mountain 4
3872 Moura 8
3873 Mouskouri 1
3874 Mozambique 4
3875 Mozart 1
3876 Moçambique 47
3877 Moçambiques 3
3878 Mr 8
3879 Mrs 12
3880 Msaccess.exe 1
3881 Mugabe 1
3882 Mulder 2
3883 Murcia 1
3884 Murphy 1
3885 Muscardini 1
3886 Musik 1
3887 Musiken 1
3888 Musselodlingen 1
3889 Mussolinihaka 1
3890 Mweta 18
3891 Mwetas 4
3892 Myanmar 2
3893 Mycket 15
3894 Myller 1
3895 Myndigheten 2
3896 Myndighetens 2
3897 Män 1
3898 Mängden 1
3899 Mängdfunktionerna 1
3900 Människor 5
3901 Människorna 4
3902 Människors 2
3903 Människorättsorganisationen 1
3904 Människorättsorganisationer 1
3905 Människorättspolitiken 1
3906 Mänskliga 9
3907 Mänsklighetens 1
3908 Märkligt 2
3909 Märks 1
3910 Mätare 1
3911 Mätt 1
3912 Må 1
3913 Måhända 1
3914 Målarfärgen 1
3915 Målet 13
3916 Målsättningen 3
3917 Många 36
3918 Månljuset 1
3919 Måste 3
3920 Måtte 2
3921 Méndez 1
3922 Möblerna 1
3923 Möjligen 1
3924 Möjligheten 3
3925 Möjligheter 1
3926 Möjligt 1
3927 Mörkt 1
3928 Möten 1
3929 München 3
3930 Münchens 1
3931 Münchhausen 1
3932 NGL-gruppen 3
3933 NL 7
3934 Nagorno-Karabach 2
3935 Namibia 6
3936 Namnet 3
3937 Namnge 1
3938 Nana 1
3939 Napoleonkrigen 1
3940 Napolitano 6
3941 Napolitanos 1
3942 Narkotikafrågan 1
3943 Narkotikahandeln 1
3944 Nasdaq 2
3945 Nasdaq- 1
3946 Nassau 3
3947 Nassaumötets 1
3948 Nasser 3
3949 Nassers 3
3950 National 2
3951 Nationaliteter 1
3952 Nationalstaterna 1
3953 Nationella 5
3954 Nationernas 4
3955 Nations 1
3956 Nato 38
3957 Nato-församlingens 1
3958 Nato-länderna 1
3959 Nato-styrkornas 1
3960 Natoaktionen 1
3961 Natobasen 1
3962 Natos 35
3963 Natostyrkor 1
3964 Natostyrkornas 1
3965 Natten 1
3966 Natura 5
3967 Naturliga 1
3968 Naturligtvis 37
3969 Neapel 2
3970 Nederländerna 25
3971 Nederländernas 1
3972 Nedläggningen 1
3973 Neil 9
3974 Neils 2
3975 Nej 32
3976 Nellie 1
3977 Ner 1
3978 Nere 1
3979 Nervcentrum 1
3980 Netanyahus 1
3981 New 15
3982 Newcastle 1
3983 News 2
3984 Newton 1
3985 Ni 176
3986 Ni-vet-vem 1
3987 Nicaragua 1
3988 Nice 1
3989 Nicholson 1
3990 Nicole 4
3991 Nicosia 1
3992 Nicosias 2
3993 Nielsen 2
3994 Nielsens 1
3995 Nielson 23
3996 Nielsons 3
3997 Nigeria 3
3998 Nikitin 2
3999 Nimbus 1
4000 Nissan 1
4001 Nivån 2
4002 Nja 1
4003 Njaa 1
4004 Nobelpris 1
4005 Nobelpristagare 1
4006 Nog 1
4007 Noggrann 1
4008 Nogueira 4
4009 Noirmoutier 1
4010 Noiz 1
4011 Nord 4
4012 Nord-Pas-de-Calais 1
4013 Nord-Syd 1
4014 Nordafrika 3
4015 Nordatlanten 2
4016 Nordatlantiska 1
4017 Norden 1
4018 Nordeuropa 1
4019 Nordirland 10
4020 Nordirlands 3
4021 Nordisk 7
4022 Norditalien 1
4023 Nordostatlantpakten 1
4024 Nordpolen 1
4025 Nordsjön 3
4026 Nordsjöområdet 1
4027 Norge 13
4028 Norges 1
4029 Normala 1
4030 Normer 1
4031 Norr 1
4032 North 1
4033 Northfield 1
4034 Now 2
4035 Now-projektet 1
4036 Noël 1
4037 Nu 74
4038 Null-värde 1
4039 Null-värden 1
4040 Null-värdet 1
4041 Numera 2
4042 Nuova 1
4043 Nuts 1
4044 Nuvarande 1
4045 Nya 8
4046 Nyckeln 1
4047 Nyexploaterade 1
4048 Nyheterna 1
4049 Nyligen 2
4050 Nyss 1
4051 Nytt 2
4052 Nyttan 2
4053 Nyttofordon 1
4054 Nz 2
4055 Nämnda 1
4056 När 330
4057 Nära 1
4058 Näringslivet 1
4059 Närmare 1
4060 Nästa 83
4061 Nästan 3
4062 Nå 3
4063 Någon 12
4064 Någonstans 1
4065 Någonting 4
4066 Något 11
4067 Några 16
4068 Nåja 3
4069 Nån 1
4070 Nåväl 3
4071 Nödvändigheten 1
4072 Nödvändigt 1
4073 Núñez 1
4074 O 1
4075 OAS 1
4076 OAU 2
4077 OAVHÄNGIGHETEN 1
4078 OCH 2
4079 OCHA 1
4080 OECD 2
4081 OECD-länderna 1
4082 OFSR 1
4083 OK 1
4084 OLAF 20
4085 OLAF:s 1
4086 OLE 2
4087 OLFAF 1
4088 OM 2
4089 OMRÖSTNING 9
4090 OSSE 1
4091 OSSE-observatörer 1
4092 OSSE:s 1
4093 OTC-derivat 10
4094 OTC-derivaten 3
4095 OTC-instrument 6
4096 OTC-instrumenten 1
4097 OTC-investeringar 1
4098 Oanmälda 1
4099 Oansvarighet 1
4100 Oavsett 7
4101 Oavslutad 1
4102 Oberbayern 1
4103 Oberoende 4
4104 Obnova-programmen 1
4105 Obs 1
4106 Och 279
4107 Också 12
4108 Odara 9
4109 Odaras 2
4110 Oddy 1
4111 Odysseus 1
4112 Offentliga 2
4113 Offentligheten 1
4114 Office 25
4115 Office-pivottabellkomponent 1
4116 Office-program 1
4117 Offret 1
4118 Ofta 3
4119 Oförfärat 1
4120 Oförmögna 1
4121 Oil 3
4122 Oil-programmet 1
4123 Ojala 1
4124 Ojeda 1
4125 Oklahoma 1
4126 Olika 3
4127 Olivia 6
4128 Olivias 1
4129 Olivier 1
4130 Oljebälte 1
4131 Oljebältet 1
4132 Oljestället 1
4133 Oljetankern 1
4134 Oljeutsläppet 1
4135 Olle 4
4136 Olyckan 2
4137 Olyckligtvis 1
4138 Olympe 1
4139 Olympic 1
4140 Om 382
4141 Omagh 1
4142 Omfånget 1
4143 Omkring 1
4144 Omlastningar 1
4145 Omorganisation 1
4146 Omräknat 1
4147 Området 3
4148 Omröstningen 56
4149 Omstrukturering 2
4150 Omstruktureringen 1
4151 Omständigheterna 1
4152 Omyndiga 1
4153 Onesta 1
4154 Online 1
4155 Onödigt 1
4156 Oomen-Ruijten 1
4157 Oostlander 3
4158 Operators 1
4159 Opinionsnätverk 1
4160 Oraninvånarnas 1
4161 Ord 3
4162 Orden 2
4163 Order 1
4164 Orderdetaljer 1
4165 Orderingången 1
4166 Ordet 6
4167 Ordförande 9
4168 Ordföranden 2
4169 Ordförandeskap 1
4170 Ordförandeskapet 9
4171 Ordförandeskapets 2
4172 Organet 1
4173 Organisationen 2
4174 Organization 1
4175 Orienten 2
4176 Orkanen 2
4177 Orkney 1
4178 Ormen 1
4179 Oron 2
4180 Oroväckande 1
4181 Orsaken 6
4182 Orsakerna 1
4183 Ortega 4
4184 Orwell 2
4185 Osip 1
4186 Oslo 3
4187 Osloavtalen 2
4188 Osloprotokollet 1
4189 Osman 1
4190 Ospar 6
4191 Ospar-avtalen 1
4192 Ospar-konventionen 3
4193 Ospar-målen 2
4194 Ospar-målet 1
4195 Ospar-normen 1
4196 Ospar-värdet 1
4197 Ostindiska 1
4198 Osäkerhet 1
4199 Otaliga 1
4200 Otroligt 1
4201 Oturligt 1
4202 Otvivelaktigt 1
4203 Ouvrière 1
4204 Oz 3
4205 PATH 1
4206 PNV 1
4207 PPE 5
4208 PPE-DE 6
4209 PPE-DE- 2
4210 PPE-DE-gruppen 3
4211 PPE-DE-gruppens 2
4212 PPE-DE-ledamöter 1
4213 PPE-gruppen 4
4214 PPE-gruppens 1
4215 PR-effekt 1
4216 PR-experter 1
4217 PR-firmor 1
4218 PSE 2
4219 PSE-gruppen 5
4220 PSE-gruppens 3
4221 PT 27
4222 PVC 3
4223 PVC-leksaker 1
4224 Pack 3
4225 Package 1
4226 Packs 2
4227 Padanien 2
4228 Paddington 2
4229 Page 2
4230 Pakistan 4
4231 Pakistans 1
4232 Palacio 18
4233 Palacios 2
4234 Palermo 1
4235 Palestina 10
4236 Palestina-Israel 1
4237 Palestinaflyktingarnas 1
4238 Palestinafrågan 1
4239 Palestinas 1
4240 Palestinierna 1
4241 Panama 1
4242 Panza 1
4243 Paolo 1
4244 Papandreou 1
4245 Papayannakis 3
4246 Papoutsis 1
4247 Pappa 2
4248 Paradoxalt 2
4249 Paragrafrytteriet 1
4250 Parallella 1
4251 Parallellt 2
4252 Paris 6
4253 Parisfördragen 1
4254 Parisprotokollet 1
4255 Park 3
4256 Parken 1
4257 Parker 1
4258 Parlament 2
4259 Parlamentet 94
4260 Parlamentets 7
4261 Parlamentsledamöterna 1
4262 Parlamentsledamöternas 1
4263 Parlement 1
4264 Partido 1
4265 Partnerskap 1
4266 Partnerskapet 1
4267 Partnerskapets 1
4268 Pas 1
4269 Passagerarna 1
4270 Patricia 1
4271 Patten 55
4272 Pattens 8
4273 Paul 6
4274 Paul-Marie 1
4275 Pays 1
4276 Pays-de-Loire 1
4277 Peake 2
4278 Pecunia 1
4279 Peijs 2
4280 Peking 2
4281 Pekingdeklarationen 1
4282 Pekingkonferensen 1
4283 Pen 1
4284 Pensioner 1
4285 Pensionsfonder 1
4286 Pensionärerna 1
4287 Pensionärspartiet 3
4288 Pentagon 1
4289 Percy 4
4290 Peres 1
4291 Perfomance 1
4292 Personalsystemet 1
4293 Personer 1
4294 Personligen 8
4295 Peter 10
4296 Peters 2
4297 Petersberg 2
4298 Petersberguppgifter 1
4299 Petersberguppgifterna 3
4300 Petersen 1
4301 Petroleum 1
4302 Pettigrew 3
4303 Pettigrews 2
4304 Petunia 9
4305 Petunias 1
4306 Phare 6
4307 Phare- 1
4308 Phare-programmen 1
4309 Phare-programmet 2
4310 Philippe 1
4311 Philoxenia-programmet 2
4312 Phonograms 1
4313 Piecyk 4
4314 Pietrasanta 1
4315 Pietro 9
4316 Pietro-betänkandet 1
4317 Pietros 4
4318 Pinochet 10
4319 Pinochet-Ugarte 1
4320 Pintassilgobetänkandet 1
4321 Piqué 1
4322 Pirker 1
4323 Pivotabellvyns 1
4324 Pivotdiagramvy 1
4325 Pivottabeller 2
4326 Pivottabellista 1
4327 Pivottabellvy 1
4328 Pjoska 1
4329 Plaid 1
4330 Planeringskommittén 1
4331 Planerna 1
4332 Plantation 1
4333 Plantin 1
4334 Plast- 1
4335 Plastindustrin 1
4336 Platons 1
4337 Plooij-van 3
4338 Plumb 1
4339 Plumb-Delors-avtalet 1
4340 Pläderingen 1
4341 Plötsligt 2
4342 Poettering 11
4343 Poetterings 1
4344 Pohjamo 1
4345 Pojkaktig 1
4346 Pojkarna 1
4347 Pojken 4
4348 Polen 6
4349 Polens 1
4350 Polisen 2
4351 Poliser 1
4352 Polisstyrkan 1
4353 Political 1
4354 Politik 1
4355 Politiken 3
4356 Politikens 1
4357 Polje 1
4358 Pollution 3
4359 Polo 1
4360 Pomés 1
4361 Ponnambalam 1
4362 Poos 4
4363 Popo 1
4364 Popular 1
4365 Port 3
4366 Portugal 36
4367 Portugals 7
4368 Portuguesa 1
4369 Positiv 1
4370 Posselt 5
4371 Post 1
4372 Post-Europa 1
4373 Posten 4
4374 Postföretaget 1
4375 Postkontoren 1
4376 Postkontorets 1
4377 Postmarknaden 1
4378 Posts 1
4379 Postsektorn 2
4380 Posttjänsten 5
4381 Posttjänster 1
4382 Posttjänsterna 5
4383 Postverken 1
4384 Potentiella 1
4385 Pottaskan 1
4386 Potter 2
4387 Poul 1
4388 Poulenc 1
4389 Power 4
4390 Prag 1
4391 Praktiskt 1
4392 Precis 17
4393 Premiärminister 1
4394 Premiärministrar 1
4395 Premiärministrarna 1
4396 Presentationen 1
4397 President 2
4398 Pressfrihet 2
4399 Presumtivt 1
4400 Preussag 1
4401 Principen 6
4402 Principförklaringar 1
4403 Prioriteringen 1
4404 Privatisering 1
4405 Privet 3
4406 Problem 2
4407 Problemen 3
4408 Problemet 19
4409 Procacci 2
4410 Procaccis 1
4411 Procentsatserna 1
4412 Processen 7
4413 Processer 1
4414 Processerna 1
4415 Prodi 103
4416 Prodi-dokument 1
4417 Prodi-kommissionen 1
4418 Prodikommissionen 1
4419 Prodis 26
4420 Producenten 1
4421 Producenternas 1
4422 Produkter 1
4423 Programmappen 1
4424 Programmen 3
4425 Programmet 7
4426 Projekt 1
4427 Projekten 2
4428 Projektet 1
4429 Prokollet 1
4430 Pronk 3
4431 Propaganda 1
4432 Property 2
4433 Protection 2
4434 Protocol 1
4435 Protokoll 1
4436 Protokollen 1
4437 Protokollet 14
4438 Provan 2
4439 Provans 1
4440 Príncipes 1
4441 Pröva 1
4442 Puerta 2
4443 Punkt 4
4444 Purvis 4
4445 Putin 2
4446 Putins 1
4447 Pyrenéerna 1
4448 PÅ 1
4449 På 163
4450 Påståendet 1
4451 Pétain 1
4452 Pöbelvälde 1
4453 QE2 1
4454 QE2:s 1
4455 Quecedo 3
4456 Queiro 1
4457 Queiró 1
4458 Quentin 1
4459 Quijote 9
4460 Quinn 85
4461 Quinns 1
4462 Quousque 1
4463 RC 1
4464 REP 2
4465 REVOKE 1
4466 RINA 3
4467 ROWS 1
4468 RSPB 1
4469 Ra-Ra 1
4470 Rabingruppen 1
4471 Racan 1
4472 Rachidi 1
4473 Rack 2
4474 Radio 4
4475 Radwan 4
4476 Rafael 4
4477 Rambeslutet 1
4478 Rambouillet 1
4479 Ramdirektivet 2
4480 Ramen 1
4481 Ramprogrammet 1
4482 Ramvillkoren 2
4483 Randzio-Plath 4
4484 Randzio-Plaths 1
4485 Raninsy 1
4486 Rapkay 8
4487 Rapkaybetänkandet 1
4488 Rapkays 2
4489 Rapporten 4
4490 Ras 3
4491 Raschhofer 1
4492 Rasismen 1
4493 Rasistiska 2
4494 Ratificeringen 1
4495 Rato 1
4496 Rauf 2
4497 Ravenna 1
4498 Rayburnspis 1
4499 Raymond 1
4500 Reactor 1
4501 Reading 1
4502 Reaktionen 1
4503 Real 1
4504 Rebecca 4
4505 Rechar-programmet 1
4506 Redan 12
4507 Redarna 1
4508 Rederiet 1
4509 Reding 7
4510 Redings 2
4511 RefLibPaths-nyckel 2
4512 Referenser 2
4513 Reformen 6
4514 Reformering 1
4515 Reformeringen 1
4516 Reformerna 1
4517 Reformprocessen 2
4518 Regensburg 1
4519 Regeringarna 1
4520 Regeringen 6
4521 Regeringsförhandlingar 1
4522 Regeringskonferensen 2
4523 Regeringskonferensens 1
4524 Regionala 1
4525 Regionalpolitiken 1
4526 Regionen 2
4527 Regioner 1
4528 Regionerna 1
4529 Regionkommittén 2
4530 Regis 1
4531 Regler 2
4532 Regleringen 1
4533 Reglerna 1
4534 Reith 1
4535 Rekommendation 1
4536 Rektorn 1
4537 Relevant 1
4538 Religionen 1
4539 Remington 1
4540 Rengie 2
4541 Rengies 1
4542 Rent 2
4543 Report 1
4544 ReportML 5
4545 ReportML-filen 1
4546 ReportML-format 1
4547 Representantgrupperna 1
4548 Republikaner 1
4549 Republiken 12
4550 Reserves 1
4551 Resolution 1
4552 Resolutionen 1
4553 Resolutionens 1
4554 Resolutioner 1
4555 Resolutionsförslag 4
4556 Resolutionsförslaget 1
4557 Resource 1
4558 Restaurant 1
4559 Resten 2
4560 Resterande 1
4561 Resterna 2
4562 Restore 1
4563 Resultat 2
4564 Resultaten 3
4565 Resultatet 9
4566 Resurser 1
4567 Retroaktiv 1
4568 Revideringen 1
4569 Revisionsrätten 5
4570 Rezala 2
4571 Rhen 1
4572 Rhendalen 1
4573 Rhenguld 2
4574 Rhenlandets 1
4575 Rhino 5
4576 Rhodesia 3
4577 Rhodesierna 1
4578 Rhone-Poulenc 1
4579 Rhône-Alpes 1
4580 Ricardo 1
4581 Richard 1
4582 Richterskalan 2
4583 Ries 1
4584 Rights 2
4585 Riis-Jørgensen 2
4586 Rika 1
4587 Riktlinjer 1
4588 Riktlinjerna 3
4589 Ringen 1
4590 Ringholm 2
4591 Rio 4
4592 Rio- 1
4593 Rio-konferensen 1
4594 Rioförklaringen 1
4595 Risken 3
4596 Ritt 1
4597 Riverside 5
4598 Road 2
4599 Robert 2
4600 Robertson 1
4601 Rocard 1
4602 Rocards 1
4603 Roissys 1
4604 Rojos 1
4605 Roland 1
4606 Rollen 2
4607 Roly 2
4608 Rom 7
4609 Rom- 1
4610 Romano 10
4611 Romfördraget 3
4612 Romfördragets 1
4613 Romkonferensen 1
4614 Romkonventionerna 1
4615 Román 2
4616 Ron 25
4617 Rons 3
4618 Roo 1
4619 Roosevelt 1
4620 Ropet 1
4621 Rosenberg 1
4622 Roth-Behrendt 10
4623 Roth-Behrendts 1
4624 Rothe 2
4625 Rotterdam 3
4626 Round 2
4627 Roure 1
4628 Rover 2
4629 Royal 2
4630 Rugby 1
4631 Rugovas 1
4632 Ruiz 1
4633 Rummet 1
4634 Rumänerna 1
4635 Rumänien 18
4636 Runt 3
4637 Rush 1
4638 Rusjailo 1
4639 Rwanda 1
4640 Ryska 1
4641 Ryssarna 1
4642 Ryssland 19
4643 Rysslands 5
4644 Räcker 1
4645 Räkna 1
4646 Rätten 1
4647 Rättsstaten 1
4648 Rättssäkerheten 1
4649 Rättstillämpningen 1
4650 Rättvisa 2
4651 Råder 1
4652 Rådet 35
4653 Rådets 17
4654 Rådsmötet 1
4655 Rådsordföranden 1
4656 Rådsordförandeskapet 1
4657 Réunion 3
4658 Röda 2
4659 Rörande 3
4660 Rösta 1
4661 Rösterna 1
4662 Röstförklaringar 1
4663 Röstförklaringar- 1
4664 Rött 1
4665 Rübig 2
4666 Rübigs 1
4667 SAP 1
4668 SCRS 1
4669 SCRS-undersökningen 1
4670 SEK 1
4671 SEK(1998 3
4672 SEK(1999)1279 2
4673 SEK(99)0066 1
4674 SELECT 1
4675 SEM-2000 1
4676 SMAKAR 1
4677 SN 1
4678 SOLAS 1
4679 SPÖ 3
4680 SQL 8
4681 SQL-fråga 1
4682 SQL-frågeläge 11
4683 SQL-frågelägen 5
4684 SQL-frågelägena 1
4685 SQL-frågeläget 1
4686 SQL-frågor 1
4687 SQL-specifikationen 1
4688 SQL-syntax 1
4689 SQL-syntaxen 1
4690 SQL-uttryck 2
4691 SQL-uttrycken 1
4692 SS 1
4693 STOA 1
4694 SUD 1
4695 SUM-DISTINCT-Pris 1
4696 Sa 1
4697 Sacharovpriset 1
4698 Sages- 1
4699 Sagorna 1
4700 Sahara 4
4701 Sahel 1
4702 Saint-Exupérys 1
4703 Saint-Josse 1
4704 Sakellariou 1
4705 Sakellarious 1
4706 Saken 1
4707 Saker 2
4708 Salafranca 2
4709 Salafrancas 1
4710 Sam 4
4711 Samarbete 3
4712 Samarbetet 2
4713 Samarbetsavtalet 1
4714 Samband 1
4715 Sambandet 1
4716 Samhällena 1
4717 Samhället 2
4718 Samma 9
4719 Sammanfattningsvis 5
4720 Sammanflätningen 1
4721 Sammanhängande 1
4722 Sammanhållningen 1
4723 Sammanhållningsfonden 15
4724 Sammanhållningsfondens 1
4725 Sammansättningen 1
4726 Sammantaget 1
4727 Sammanträdena 1
4728 Sammanträdet 23
4729 Samordning 3
4730 Samordningen 1
4731 Samstämmighet 1
4732 Samstämmigheten 3
4733 Samtal 1
4734 Samtalen 1
4735 Samtidigt 43
4736 Samtliga 5
4737 San 2
4738 Sancho 1
4739 Sandbankar 1
4740 Sandbæk 1
4741 Sanningen 8
4742 Sanningens 1
4743 Sannolikt 1
4744 Santa 1
4745 Santer 3
4746 Santer-kommissionen 1
4747 Santer-kommissionens 1
4748 Santerkommissionens 1
4749 Santiago 1
4750 Santos 3
4751 Sapar 1
4752 Sapard 3
4753 Saramago 2
4754 Sardinernas 1
4755 Sarre-Lorraine-Luxemburg 1
4756 Saudiarabien 1
4757 Save 6
4758 Save- 1
4759 Save-programmet 2
4760 Savefloden 1
4761 Savimbi 1
4762 Savimbis 1
4763 Scarborough 1
4764 Scenen 1
4765 Scharping 1
4766 Scheele 1
4767 Schengen 3
4768 Schengenavtalen 1
4769 Schengenavtalet 3
4770 Schengenkonventionen 1
4771 Schengenkonventionens 1
4772 Schengenområdet 1
4773 Schengenregelverket 1
4774 Schengenstat 1
4775 Schierhuber 1
4776 Schipol-flygplats 1
4777 Schleicher 3
4778 Schmid 1
4779 Schmidbetänkandet 1
4780 Schmidt 10
4781 Schmidtbetänkandet 1
4782 Schmidts 4
4783 Schori 2
4784 Schreyer 4
4785 Schroedter 10
4786 Schroedterbetänkandet 2
4787 Schroedters 6
4788 Schröder 1
4789 Schultz 2
4790 Schulz 7
4791 Schwaigerbetänkandet 1
4792 Schwarzwald 1
4793 Schweiz 3
4794 Schörling 1
4795 Schüssel 6
4796 Schüssels 1
4797 Sdot 1
4798 Se 5
4799 Sea 1
4800 Seattle 23
4801 Sebastian 1
4802 Sedan 67
4803 Sedvänjorna 1
4804 Segni 1
4805 Segura 1
4806 Seguro 1
4807 Seixas 6
4808 Sekelgammal 1
4809 Sektorn 1
4810 Sellafield 1
4811 Seminarier 1
4812 Sen 7
4813 Senare 3
4814 Senast 1
4815 Sens 1
4816 Sent 1
4817 Seppänen 1
4818 Ser 1
4819 Serbien 32
4820 Serbiens 4
4821 Seriösa 1
4822 Server-databas 1
4823 Service 1
4824 Sett 1
4825 Sevilla 1
4826 Sex 3
4827 Sha'ananim 1
4828 Shahar 5
4829 Shaping 3
4830 Sharm 4
4831 Sharm-el-Sheik 1
4832 Shell 3
4833 Shepherdstown 3
4834 Shetland 1
4835 Shetlandsöarna 2
4836 Shimon 1
4837 Shinza 3
4838 Shinzas 1
4839 Shipping 2
4840 Shop 1
4841 Short 1
4842 Sibirien 1
4843 Sicilien 1
4844 Siciliens 1
4845 Sid 1
4846 Side 1
4847 Sidor 1
4848 Siena 1
4849 Sierra 1
4850 Sifferuppgifterna 1
4851 Siffran 1
4852 Siffrorna 1
4853 Sihanouk 1
4854 Sikten 1
4855 Silver 4
4856 Simpson 1
4857 Sin 1
4858 Sinjavskij 2
4859 Sintra 8
4860 Sintraavtal 1
4861 Sintrafördraget 1
4862 Sions 1
4863 Siri 2
4864 Sist 2
4865 Sisyfosarbete 1
4866 Sisyfosklippa 1
4867 Situationen 15
4868 Sju 1
4869 Sjukdomen 3
4870 Sjukhusläkare 1
4871 Sjukvård 1
4872 Själv 5
4873 Själva 4
4874 Självfallet 1
4875 Självklart 5
4876 Sjätte 2
4877 Sjömäns 1
4878 Sjöstedt 7
4879 Sjötransporten 1
4880 Ska 3
4881 Skadestånd 1
4882 Skador 1
4883 Skadorna 1
4884 Skall 9
4885 Skapa 1
4886 Skapandet 3
4887 Skaror 1
4888 Skattedebiteringen 1
4889 Skatteharmonisering 1
4890 Skeppet 1
4891 Sker 1
4892 Skillnaderna 3
4893 Skjulet 1
4894 Skogsvårdsmyndigheten 1
4895 Skopje 4
4896 Skotsk 1
4897 Skottland 25
4898 Skottlands 2
4899 Skrapie 1
4900 Skulden 1
4901 Skulle 22
4902 Skvallret 1
4903 Skydd 2
4904 Skyddet 4
4905 Skyddsåtgärderna 1
4906 Skyltar 1
4907 Skälen 1
4908 Skälet 6
4909 Slapphet 1
4910 Slovakien 1
4911 Slovenien 1
4912 Slut 1
4913 Sluta 1
4914 Slutligen 82
4915 Slutrapporten 1
4916 Slutresultatet 2
4917 Slutsatsen 3
4918 Slutsatserna 4
4919 Släpp 1
4920 Släppområden 3
4921 Släppområdena 1
4922 Smith 2
4923 Smiths 1
4924 Små 1
4925 Småföretagare 1
4926 Snabb 1
4927 Snarare 3
4928 Snart 1
4929 Snödrottningsspegel 1
4930 Soares 3
4931 Social 1
4932 Socialfonden 2
4933 Socialistgruppen 1
4934 Socialpolitik 1
4935 Socialpolitiken 2
4936 Socialpolitiska 1
4937 Society 1
4938 Soekarnopoetri 1
4939 Sokrates- 1
4940 Solana 52
4941 Solanas 4
4942 Solbes 6
4943 Soldat 1
4944 Soldater 1
4945 Solen 5
4946 Solidaritet 1
4947 Solidariteten 1
4948 Solsjenitsyns 1
4949 Som 180
4950 Somalia 1
4951 Somes 2
4952 Somliga 7
4953 Souchet 2
4954 Souladakis 2
4955 Southampton 2
4956 Souto 1
4957 Sovjetunionen 2
4958 Sovjetunionens 1
4959 Spanien 52
4960 Spaniens 4
4961 Spara 5
4962 Spararna 1
4963 Speciella 1
4964 Speciellt 1
4965 Specifika 2
4966 Spegelbilden 1
4967 Spelar 1
4968 Spencer 1
4969 Speroni 1
4970 Spindlarna 1
4971 Sport 1
4972 Spridda 1
4973 Språket 1
4974 Sputnikbaren 5
4975 Sr 1
4976 Sri 3
4977 St 5
4978 Stabex- 1
4979 Stabiliserings- 1
4980 Stabiliteten 1
4981 Stabilitetspakten 3
4982 Stabilitetspaktens 1
4983 Stackars 4
4984 Staden 1
4985 Stadens 1
4986 Stadgan 3
4987 Stadsmiljöpolitiken 1
4988 Staes 1
4989 Stafford 1
4990 Standardinställningen 1
4991 Standardläge 1
4992 Standardläget 1
4993 Stanna 1
4994 Start- 1
4995 Stater 1
4996 Staterna 6
4997 Staternas 1
4998 Stationerna 1
4999 Statistiken 1
5000 Statlig 1
5001 Statliga 2
5002 Statligt 1
5003 Statsbalen 1
5004 Statsmakten 1
5005 Steel 1
5006 Stegrennan 1
5007 Stegrennans 3
5008 Stegrennansstrandremsa 1
5009 Stella 5
5010 Stenar 1
5011 Stendhals 1
5012 Stenmarck 2
5013 Stenzel 8
5014 Stenzels 6
5015 Stephen 2
5016 Sterckx 5
5017 Stickordet 1
5018 Stilla 4
5019 Stillahavsområdet 2
5020 Stillman 44
5021 Stillmans 8
5022 Stockholm 5
5023 Stoke-on-Trent 1
5024 Stolarna 1
5025 Stora 4
5026 Storbritannien 25
5027 Storbritanniens 2
5028 Storebror 1
5029 Storhertigdömet 1
5030 Stormar 1
5031 Stormarna 1
5032 Stormen 1
5033 Storskalig 1
5034 Stort 1
5035 Straffrätten 1
5036 Straffrättslig 1
5037 Straffrättsliga 1
5038 Straffångar 1
5039 Strasbourg 26
5040 Strasbourgförklaringen 2
5041 Strasbourgs 1
5042 Strategidokumentet 1
5043 Strategiska 1
5044 Stravinskij 1
5045 Strax 1
5046 Street 2
5047 Stregrennan 1
5048 Stromboli 2
5049 Strukturellt 2
5050 Strukturfonderna 2
5051 Strukturfondernas 2
5052 Sträng 1
5053 Strävan 1
5054 Strävar 1
5055 Strålande 1
5056 Strömmen 1
5057 Studenter 1
5058 Studies 1
5059 Style 1
5060 Stylesheet 2
5061 Styrkan 1
5062 Städerna 1
5063 Stämmer 2
5064 Stämningen 1
5065 Ständiga 1
5066 Stålsektorn 1
5067 Ståndpunkterna 1
5068 Står 1
5069 Stöd 5
5070 Stöden 1
5071 Stöder 2
5072 Stödpunkten 1
5073 Stödsystemet 1
5074 Större 2
5075 Största 2
5076 Suanzes-Carpegna 4
5077 Subsidiariteten 1
5078 Subventioner 2
5079 Suckande 1
5080 Sudan 3
5081 Sudre 2
5082 Suffolk 1
5083 Sui 1
5084 Suisse 1
5085 Summan 1
5086 Suominen 2
5087 Suveräniteten 1
5088 Svaret 5
5089 Svart 1
5090 Svarta 1
5091 Svartvändargränden 2
5092 Svend 1
5093 Svenska 2
5094 Svepeskålen 1
5095 Sverige 44
5096 Sveriges 3
5097 Svårigheten 3
5098 Svårigheterna 1
5099 Swaziland 2
5100 Swoboda 15
5101 Swobodabetänkandet 1
5102 Swobodas 7
5103 Syd 8
5104 Sydafrika 22
5105 Sydafrikaavtalen 1
5106 Sydafrikas 2
5107 Sydamerika 2
5108 Sydeuropa 3
5109 Sydkorea 1
5110 Sydostasien 3
5111 Sydosteuropa 1
5112 Sydösteuropa 2
5113 Syftet 20
5114 Synd 1
5115 Synnerligen 1
5116 Syrien 26
5117 Syriens 2
5118 Syrierna 2
5119 Sysminsystemet 1
5120 Sysselsättningen 4
5121 Sysselsättningspakten 1
5122 Sysselsättningsstrategin 1
5123 System 1
5124 System32 1
5125 Systemen 1
5126 Systemmappen 1
5127 Sánchez 3
5128 São 2
5129 Säg 2
5130 Säger 1
5131 Säker 1
5132 Säkerheten 1
5133 Säkerhetsaspekten 1
5134 Säkerhetskoefficienten 1
5135 Säkerhetsrådgivare 1
5136 Säkerhetsåtgärderna 1
5137 Säkerligen 2
5138 Säkert 1
5139 Sämre 1
5140 Särskild 2
5141 Särskilda 1
5142 Särskilt 12
5143 Säsongen 1
5144 Sättet 1
5145 Så 95
5146 Sådan 2
5147 Sådana 16
5148 Sådant 1
5149 Således 14
5150 Sålunda 3
5151 Såna 1
5152 Sången 1
5153 Sånt 2
5154 Såsom 9
5155 Såvitt 3
5156 Såväl 6
5157 Sète 1
5158 Söder 1
5159 Söderhavet 1
5160 Söderman 1
5161 Södermans 1
5162 Södern 1
5163 Sökvägarna 1
5164 Sörensen 1
5165 T-tack 1
5166 T.ex. 1
5167 T.o.m. 1
5168 TBT 3
5169 TDI-gruppen 3
5170 TO 1
5171 TRIPS 1
5172 TRIPS-avtalen 2
5173 TSE 5
5174 TSE-risker 1
5175 TSE-sjukdomar 3
5176 TV 8
5177 TV-apparaten 1
5178 TV-apparater 1
5179 TV-bevakningen 1
5180 TV-bilder 1
5181 TV-bilderna 1
5182 TV-bolagen 1
5183 TV-kanal 4
5184 TV-kanalen 2
5185 TV-kanaler 3
5186 TV-program 2
5187 TV-programmen 1
5188 TV-skärmar 1
5189 TV-skärmen 1
5190 TV-sändare 1
5191 TV-team 1
5192 TV-tekniker 1
5193 TV-torn 1
5194 TV-utsändningar 1
5195 TV:n 1
5196 Ta 14
5197 Table 1
5198 Tacis 4
5199 Tacis- 1
5200 Tacis-programmet 2
5201 Tack 126
5202 Tadzjikistan 5
5203 Tag 1
5204 Taiwan 1
5205 Tajani 1
5206 Tajo-Segura- 1
5207 Tal 1
5208 Tala 2
5209 Talar 5
5210 Talaren 1
5211 Talmannen 24
5212 Tammerfors 33
5213 Tammerforsavtalen 1
5214 Tammerforsbeslutens 1
5215 Tang 1
5216 Tanganyika 1
5217 Tanio 1
5218 Tanken 5
5219 Tanzania 2
5220 Tar 1
5221 Tarek 1
5222 Tas 1
5223 Tauerntunneln 1
5224 Taxis 1
5225 Tecken 1
5226 Tekniska 2
5227 Telefonen 1
5228 Telekommunikationsministeriet 1
5229 Teresa 1
5230 Terror 1
5231 Terrorism 1
5232 Terroristerna 1
5233 Terrón 5
5234 Tesauro 1
5235 Texas 2
5236 Texten 3
5237 Thaci 1
5238 Thailand 1
5239 The 5
5240 Theato 12
5241 Theatobetänkandet 1
5242 Theatos 12
5243 Themsenmynningen 2
5244 Themsenvatten 1
5245 Theo 1
5246 Theonas 2
5247 Thermonuclear 1
5248 Thompson 1
5249 Thompsons 1
5250 Thors 3
5251 Thurber 1
5252 Thurn 1
5253 Thyssen 3
5254 Thyssens 2
5255 Tibet 22
5256 Tibet-frågan 1
5257 Tiden 2
5258 Tidigare 7
5259 Tidningsartiklarna 1
5260 Tidsfristen 1
5261 Tidvattnet 1
5262 Tiffanys 1
5263 Till 101
5264 Tillfälligheter 1
5265 Tillförlitliga 1
5266 Tillgänglig 1
5267 Tillgången 1
5268 Tillhörande 1
5269 Tillsammans 4
5270 Tillståndet 2
5271 Tillverkarna 2
5272 Tillverkningen 1
5273 Tillväxt 2
5274 Tillväxten 1
5275 Tillämpning 1
5276 Tillämpningen 2
5277 Tillåt 15
5278 TillåtBorttagning 1
5279 TillåtRedigering 1
5280 TillåtTillägg 1
5281 Tillåter 3
5282 Timor 4
5283 Timothy 5
5284 Tindi 2
5285 Tingesten 1
5286 Tio 2
5287 Tiotusentals 1
5288 Tisza 3
5289 Titanic 1
5290 Titley 2
5291 Titleys 1
5292 Titta 1
5293 Tja 2
5294 Tjeckien 2
5295 Tjeckiens 2
5296 Tjernobyl 1
5297 Tjetjenien 15
5298 Tjetjenienpolitik 1
5299 Tjugo 2
5300 Tjuvars 1
5301 Tjänstekvaliteten 1
5302 Tjänsternas 1
5303 Tobin-skatt 1
5304 Today 1
5305 Toddyblom 1
5306 Todinskatten 1
5307 Tokyo 1
5308 Toledo 1
5309 Tom 1
5310 Tomma 2
5311 Tomé 2
5312 Tongivande 1
5313 Tonvikten 3
5314 Tool 1
5315 Toppmötena 1
5316 Toppmötet 5
5317 Torrey 3
5318 Torry 1
5319 Torsdag 1
5320 Torv 1
5321 Torven 1
5322 Total 8
5323 Total-Elf 1
5324 Total-Fina 3
5325 TotalFina 1
5326 Tour 1
5327 Toyota 1
5328 Trade-Related 1
5329 Tradition 1
5330 Traditionen 1
5331 Traditionsmässigt 1
5332 Trafalgar 1
5333 Trafiken 1
5334 Trafiksäkerheten 1
5335 Transformation 2
5336 Transitional 1
5337 Transnationella 1
5338 Transport 1
5339 Transportsäkerheten 1
5340 Trastfältet 1
5341 Travel 1
5342 Tre 6
5343 Treaty 2
5344 Tredje 1
5345 Trentin 1
5346 Trepca 1
5347 Tretti 1
5348 Trettiotre 1
5349 Trident 2
5350 Tridentbasen 1
5351 Trittin 1
5352 Tro 1
5353 Trojkan 1
5354 Trolla 1
5355 Trollkarlar 1
5356 Tror 12
5357 Trots 44
5358 Trovärdigheten 2
5359 Trygghetsfrågor 1
5360 Träd 1
5361 Tsatsos 6
5362 Tulsa 1
5363 Tunisien 1
5364 Tupperware 1
5365 Tupperwarekvällar 1
5366 Turin 1
5367 Turism 3
5368 Turismen 8
5369 Turismens 1
5370 Turistpolitiken 1
5371 Turkiet 72
5372 Turkiets 15
5373 Turkmenistan 2
5374 Tusen 1
5375 Tusentals 1
5376 Tvillingarnas 1
5377 Tvärs 1
5378 Tvärt 2
5379 Tvärtom 13
5380 Två 17
5381 Tvåtusen 1
5382 Ty 16
5383 Tycker 2
5384 Tyckte 1
5385 Tydliga 1
5386 Tydligen 2
5387 Tydligt 1
5388 Tyskland 40
5389 Tysklands 2
5390 Tystnaden 1
5391 Tyvärr 35
5392 Tänk 12
5393 Tänker 2
5394 Tågkraschen 1
5395 U 4
5396 U-länderna 1
5397 U-ländernas 1
5398 UCITS 4
5399 UCITS-direktivet 1
5400 UCK 5
5401 UCK-ledaren 1
5402 UCK:s 2
5403 UCLAF 1
5404 UDB 2
5405 UEN 1
5406 UEN-gruppen 3
5407 UNCTAD 1
5408 UNEF 1
5409 UNHCR 1
5410 UNIFIL 1
5411 UNITA 2
5412 UNITA-flygplatserna 1
5413 UNITA:s 2
5414 UNMIK 6
5415 US-dollar 1
5416 USA 36
5417 USA:s 2
5418 USD 1
5419 Uganda 1
5420 Ugglan 1
5421 Ukraina 2
5422 Ulster 2
5423 Undantag 1
5424 Undantagen 1
5425 Undantaget 1
5426 Under 108
5427 Underbart 1
5428 Underformulär 2
5429 Underlaget 1
5430 Underpunkten 1
5431 Undersökningarna 1
5432 Unga 1
5433 Ungdoms- 1
5434 Ungefär 2
5435 Ungern 6
5436 Ungerns 1
5437 Unice 2
5438 Unicef 1
5439 Unilever 1
5440 Union 2
5441 Unionen 24
5442 Unionens 5
5443 United 1
5444 Universal 1
5445 Universum 1
5446 Uppassare 1
5447 Uppbyggnaden 1
5448 Uppdateringen 1
5449 Uppenbarligen 3
5450 Uppfylls 1
5451 Uppföljning 2
5452 Uppgiften 3
5453 Uppgiftslämnare 1
5454 Uppgörelsen 1
5455 Upphovsmannarättigheter 1
5456 Upphovsrättsinnehavare 1
5457 Uppriktigt 2
5458 Upprättandet 2
5459 Uppsikt 1
5460 Ur 19
5461 Urba- 1
5462 Urban 27
5463 Urban-betänkandet 1
5464 Urban-dagordning 1
5465 Urban-initiativ 1
5466 Urban-initiativet 6
5467 Urban-initiativets 1
5468 Urban-program 1
5469 Urban-programmen 1
5470 Urban-programmet 12
5471 Urban-projekten 4
5472 Urban-utvecklingspolitik 1
5473 Urbans 1
5474 Urquiola 2
5475 Ursprungligen 1
5476 Ursprungsbefolkningen 2
5477 Ursprungstexten 1
5478 Ursula 2
5479 Ursäkta 6
5480 Uruguayrundan 2
5481 Urvalskriterierna 1
5482 Usted 1
5483 Ut 1
5484 Utan 20
5485 Utanför 3
5486 Utarbetandet 1
5487 Utarmningen 1
5488 Utbildning 1
5489 Utbildningen 1
5490 Utbildningsministeriet 1
5491 Utdelningen 1
5492 Utestående 1
5493 Utflödet 1
5494 Utformningen 3
5495 Utförande 1
5496 Utgiften 1
5497 Utgifterna 1
5498 Utifrån 5
5499 Utkastet 2
5500 Utmaningarna 1
5501 Utmaningen 3
5502 Utmärkt 3
5503 Utnyttjandet 1
5504 Utnämning 1
5505 Utnämningen 1
5506 Utom 1
5507 Utskottet 24
5508 Utskottets 1
5509 Utsläppet 1
5510 Uttalande 1
5511 Uttalandena 1
5512 Uttjänta 1
5513 Uttryck 1
5514 Utvecklandet 1
5515 Utvecklaren 1
5516 Utvecklingen 5
5517 Utvecklingsländer 1
5518 Utvecklingspartnerskapen 2
5519 Utvecklingssamarbetets 1
5520 Utvidgning 2
5521 Utvidgningen 5
5522 Utvidgningens 1
5523 Utvärdera 1
5524 Utöver 3
5525 Uzbekistan 2
5526 V 7
5527 V-ställda 1
5528 V. 1
5529 VBA 1
5530 VD 1
5531 VEU 5
5532 VI 2
5533 VIII 2
5534 Vaclav 6
5535 Vad 247
5536 Vadan 1
5537 Valdez 1
5538 Valdez-katastrofen 2
5539 Valen 1
5540 Valencias 1
5541 Valentins 1
5542 Valet 2
5543 Valette 1
5544 Valle 1
5545 Vallelersundi 4
5546 Vallonien 1
5547 Valverdes 1
5548 Van 15
5549 Vandamaffärerna 1
5550 Vanligen 1
5551 Vanligtvis 1
5552 Vanurå 1
5553 Vapen 1
5554 Var 24
5555 Vare 4
5556 Varela 4
5557 Varelsen 1
5558 Varenda 3
5559 Varför 54
5560 Varifrån 1
5561 Varje 37
5562 Varken 7
5563 Varning 1
5564 Varor 1
5565 Vart 3
5566 Vatanen 3
5567 Vatten 12
5568 Vattenbruket 1
5569 Vattenfrågan 1
5570 Vattenproblemet 1
5571 Vattnet 5
5572 Velzen 2
5573 Vem 24
5574 Vems 2
5575 Vendée 6
5576 Venetia 4
5577 Venezuela 2
5578 Venstres 2
5579 Ventimiglia 1
5580 Verheugen 8
5581 Verkligheten 2
5582 Verksamheten 2
5583 Verksamhetsområdet 1
5584 Verktyg-menyn 1
5585 Vermeers 1
5586 Vernon 19
5587 Vernons 4
5588 Versailles 1
5589 Verts 4
5590 Verts-gruppens 1
5591 Vet 2
5592 Vetenskapen 1
5593 Vetenskapsmännen 2
5594 Veteranbilarnas 1
5595 Vetskapen 1
5596 Vi 1650
5597 Via 4
5598 Vice 1
5599 Viceconte 6
5600 Vicecontes 4
5601 Vichyregimens 1
5602 Vid 61
5603 Vidal-Quadras 1
5604 Vidare 27
5605 Vigo 1
5606 Vikten 1
5607 Viktiga 4
5608 Viktigast 3
5609 Vilagarcia 1
5610 Vild 1
5611 Vilda 2
5612 Viljan 1
5613 Vilka 39
5614 Vilken 17
5615 Vilket 7
5616 Vill 14
5617 Ville 2
5618 Villiers 5
5619 Villkoren 2
5620 Villkorsstyrd 1
5621 Vilse 1
5622 Vin 1
5623 Vinci 2
5624 Vinden 2
5625 Vinter 1
5626 Vintergatan 3
5627 Viout 1
5628 Vireaid 1
5629 Virginia 8
5630 Viruset 2
5631 Visa 2
5632 Vissa 34
5633 Visserligen 7
5634 Visst 10
5635 Visual 3
5636 Vit 1
5637 Vita 1
5638 Vitboken 3
5639 Vitheten 1
5640 Vitoria 2
5641 Vitorino 13
5642 Vitorinos 4
5643 Vivianne 1
5644 Vivien 5
5645 Vivienne 1
5646 Vlaams 1
5647 Vlaamsblok 1
5648 Vladimir 3
5649 Vodafone-Mannesmann 1
5650 Voinet 1
5651 Vojvodina 1
5652 Voldemort 5
5653 Voldemorts 2
5654 Volksunie 1
5655 Volkswagen 1
5656 Von 1
5657 Vore 1
5658 Vraket 1
5659 Vägen 3
5660 Vägkontroller 1
5661 Väldigt 1
5662 Välj 1
5663 Väljer 2
5664 Välkommen 1
5665 Välkomsthälsning 3
5666 Vänstern 1
5667 Vänsterns 1
5668 Vänta 1
5669 Väntade 1
5670 Väntar 1
5671 Värden 1
5672 Värderade 2
5673 Världen 2
5674 Världens 1
5675 Världsbanken 4
5676 Världsbankens 1
5677 Världshandelsorganisationen 8
5678 Världshandelsorganisationens 5
5679 Världshälsoorganisationen 1
5680 Världshälsoorganisationens 2
5681 Världsnaturfonden 3
5682 Världspostföreningens 1
5683 Världssamfundet 2
5684 Värmen 1
5685 Västafrika 1
5686 Västatlantens 1
5687 Västbanken 4
5688 Västeuropa 1
5689 Västeuropeiska 3
5690 Västfrika 1
5691 Västindien 5
5692 Västmakterna 1
5693 Västprovinsen 1
5694 Västra 1
5695 Västsahara 1
5696 Västtyskland 1
5697 Västtysklands 1
5698 Växthuseffekten 1
5699 Våld 1
5700 Våldet 2
5701 Vår 55
5702 Våra 19
5703 Vårt 19
5704 Véronique 1
5705 W3C 1
5706 WCT 1
5707 WHERE 1
5708 WHO 1
5709 WINNT 1
5710 WIPO 5
5711 WIPO-avtalen 5
5712 WIPO-avtalet 10
5713 WIPO-fördragen 1
5714 WIPO-församlingen 1
5715 WIPO-överläggningar 1
5716 WIPO:s 1
5717 WPPT 1
5718 WTO 12
5719 WTO-förenlig 1
5720 WTO-förhandlingarna 1
5721 WTO-systemet 1
5722 WTO:s 5
5723 WWF 1
5724 Waddenzee 1
5725 Waffen 1
5726 Waffen-SS:s 1
5727 Wagners 1
5728 Wahid 2
5729 Wales 18
5730 Wall 1
5731 Wallström 16
5732 Wallströms 2
5733 Walter 2
5734 Warszawa 1
5735 Warszawas 1
5736 Washington 4
5737 Washingtons 3
5738 Watch 1
5739 Waterfold 1
5740 Watts 1
5741 Weasley 19
5742 Weasleys 3
5743 Web 8
5744 Webbsidans 1
5745 Weiler 1
5746 Wellington 1
5747 Wentz 18
5748 Wentz' 1
5749 West 3
5750 Westminster 1
5751 Where 1
5752 Wide 3
5753 Wiebenga 2
5754 Wieland 4
5755 Wien 4
5756 Wijkman 2
5757 Wijkmans 2
5758 Wilhelmshaven 1
5759 William 3
5760 Wilson 3
5761 Wiltshire 1
5762 Windows 2
5763 Windows-registret 1
5764 Winwardöarna 2
5765 Witness 1
5766 Wogau 18
5767 Wogaubetänkandet 1
5768 Wogaus 3
5769 Wolfsonstiftelsen 1
5770 Women 1
5771 Word 1
5772 Work 1
5773 World 7
5774 Wulf-Mathies 5
5775 Wuori 1
5776 Wurtz 10
5777 Wye 1
5778 Wye-avtalen 1
5779 Wye-avtalet 1
5780 Wynn 1
5781 X 1
5782 XI 2
5783 XML 5
5784 XML-baserade 2
5785 XML-baserat 1
5786 XML-dokument 17
5787 XML-fil 5
5788 XML-filer 2
5789 XML-informationen 2
5790 XML-källan 1
5791 XML-liknande 1
5792 XML-märken 2
5793 XML-schemafil 2
5794 XML-schemastandarden 1
5795 XML-standardformat 1
5796 XML-syntaxen 1
5797 XP 5
5798 XP-licens 5
5799 XP-licenser 1
5800 XP-nätverkslicens 1
5801 XP-program 2
5802 XSD 2
5803 XSL-fil 1
5804 XSL-formatmall 1
5805 XSL-formatmallar 1
5806 XSL-transformationsfil 1
5807 XSLT 5
5808 XX 1
5809 XXVII:e 1
5810 XXVIII:e 1
5811 Yam 1
5812 Yarmouth 1
5813 Yasser 1
5814 Yassir 1
5815 Yawlen 1
5816 Yeu 1
5817 York 11
5818 Yorker 1
5819 Yorkshire 3
5820 You 1
5821 Youngblood 1
5822 Youth 1
5823 Youthstart 2
5824 Yr 1
5825 Yrkandet 1
5826 Yrkesutbildning 1
5827 Ytterligare 3
5828 Ytterst 2
5829 Yttersta 1
5830 Yttrandet 1
5831 Yttre 3
5832 Zaire 1
5833 Zakaria 1
5834 Zambia 3
5835 Zeeland 3
5836 Zeus 8
5837 Zimbabwe 1
5838 Zimeray 1
5839 Zimmerling 1
5840 Zion 1
5841 [ 6
5842 ] 7
5843 _ 1
5844 a 19
5845 abonnentförteckningen 1
5846 absolut 126
5847 absoluta 7
5848 absorberad 1
5849 absorberade 2
5850 abstrakt 3
5851 absurd 3
5852 absurda 2
5853 absurditet 1
5854 absurt 5
5855 acceleration 1
5856 accelererande 1
5857 accentuerar 1
5858 accentueras 2
5859 accentueringarna 1
5860 acceptabel 2
5861 acceptabelt 8
5862 acceptabla 1
5863 acceptans 6
5864 acceptansen 2
5865 acceptansnivån 1
5866 acceptera 59
5867 accepterad 1
5868 accepterade 5
5869 accepterande 2
5870 accepterandet 1
5871 accepterar 18
5872 accepteras 18
5873 accepterat 7
5874 accepterats 5
5875 accountability 1
5876 ach 1
5877 ackumulerat 1
5878 acquis 3
5879 acquisition 1
5880 ad 5
5881 adderar 1
5882 additionalitet 3
5883 additionaliteten 1
5884 additionalitets- 1
5885 additionalitetsprincipen 7
5886 additionella 3
5887 adekvat 6
5888 adekvata 2
5889 adelsskap 1
5890 adjektiv 2
5891 adjektivet 1
5892 administration 8
5893 administrationen 7
5894 administrationer 1
5895 administrativ 6
5896 administrativa 29
5897 administrativt 9
5898 administratörer 1
5899 administrera 1
5900 administreras 1
5901 adriatiska 3
5902 advokat 4
5903 advokaten 1
5904 advokater 2
5905 affär 7
5906 affären 2
5907 affärer 7
5908 affärsbeslut 1
5909 affärsföretag 1
5910 affärsgrenar 1
5911 affärshemligheter 1
5912 affärslivets 1
5913 affärsmannahänder 1
5914 affärsmän 1
5915 affärsmännens 1
5916 affärsmässig 1
5917 affärspaketverksamhet 1
5918 affärsrisker 2
5919 affärsstrukturer 1
5920 affärsstrukturerna 1
5921 afrikaner 2
5922 afrikanerna 1
5923 afrikansk 1
5924 afrikanska 11
5925 afrikanskt 3
5926 aftonskolan 1
5927 age 1
5928 agenda 6
5929 agendan 3
5930 agent 2
5931 agenterna 1
5932 agera 56
5933 agerade 2
5934 agerande 42
5935 agerandet 2
5936 agerar 15
5937 agerat 6
5938 agg 1
5939 agglomerationscentra 1
5940 aggregat 1
5941 aggregaten 1
5942 aggression 3
5943 aggressioner 1
5944 aggressiv 1
5945 aggressiva 2
5946 agitation 1
5947 agrara 1
5948 agronomisk 1
5949 agroturismen 1
5950 aid 1
5951 aids 10
5952 aids-situationen 1
5953 aidsbekämpning 1
5954 aidsepidemi 1
5955 aidspatienter 2
5956 aidsrelaterad 1
5957 aidsrelaterade 1
5958 aidssiffrorna 1
5959 aidsviruset 2
5960 ajournering 2
5961 akademisk 1
5962 akademiska 1
5963 akt 18
5964 akta 3
5965 aktat 1
5966 akten 1
5967 aktens 1
5968 akter 2
5969 akterna 3
5970 akterut 1
5971 akteröver 1
5972 aktie 1
5973 aktiebolag 1
5974 aktiebolagen 1
5975 aktiebolaget 3
5976 aktiebörserna 1
5977 aktiefonder 2
5978 aktieindex 1
5979 aktieinnehav 1
5980 aktieinvesteringar 1
5981 aktiekurserna 1
5982 aktiemarknaden 2
5983 aktiemarknader 1
5984 aktier 3
5985 aktierna 2
5986 aktieägare 3
5987 aktieägarna 2
5988 aktieägarnas 2
5989 aktion 6
5990 aktionen 2
5991 aktioner 7
5992 aktionerna 3
5993 aktionsgrupper 3
5994 aktionsgrupperna 1
5995 aktionsradie 1
5996 aktiv 23
5997 aktiva 15
5998 aktivare 5
5999 aktivera 2
6000 aktiveras 3
6001 aktivering 1
6002 aktivism 1
6003 aktivistiska 1
6004 aktivitet 10
6005 aktiviteten 2
6006 aktiviteter 13
6007 aktiviteterna 4
6008 aktiviteters 1
6009 aktivitetsbaserad 1
6010 aktivitetsbaserade 1
6011 aktivt 30
6012 aktning 2
6013 aktningsbetygelse 1
6014 aktningsvärda 2
6015 aktris 1
6016 aktualisera 2
6017 aktualiseras 2
6018 aktualisering 2
6019 aktuell 9
6020 aktuella 70
6021 aktuellare 2
6022 aktuellt 8
6023 aktör 3
6024 aktören 2
6025 aktörer 27
6026 aktörerna 18
6027 aktörernas 3
6028 aktörers 2
6029 akut 6
6030 akuta 8
6031 akvarelltonade 1
6032 akvavit 3
6033 al-Sharas 1
6034 alarmerande 4
6035 alban 1
6036 albaner 7
6037 albanerna 1
6038 albansk 2
6039 albanska 13
6040 albansktalande 1
6041 aldrig 141
6042 alert 1
6043 alf 1
6044 alfabetet 1
6045 alfabetiseringsnivå 1
6046 alfer 1
6047 algbekämpning 1
6048 alias 3
6049 aliasnamn 1
6050 alibi 2
6051 alkemister 1
6052 alkohol 8
6053 alkoholbeskattning 1
6054 alkoholen 1
6055 alkoholens 1
6056 alkoholhalten 1
6057 alkoholhaltiga 7
6058 alkoholkonsumtion 1
6059 alkoholkonsumtionen 3
6060 alkoholmissbruk 1
6061 alkoholmonopol 1
6062 alkoholmonopolet 2
6063 alkoholpolitiken 2
6064 alkoholprodukter 4
6065 alkor 1
6066 all 114
6067 alla 1221
6068 allas 21
6069 alldaglig 1
6070 alldeles 95
6071 allegorisk 1
6072 allegoriska 1
6073 allehanda 4
6074 allena 1
6075 allenarådande 1
6076 allergiska 1
6077 allesammans 13
6078 allestädes 1
6079 alleuropeisk 1
6080 alleuropeiskt 2
6081 allians 5
6082 alliansen 23
6083 allianser 2
6084 alliansfria 1
6085 allierad 2
6086 allierade 3
6087 allihop 5
6088 allihopa 1
6089 allmosor 1
6090 allmän 53
6091 allmängiltiga 1
6092 allmängiltigt 1
6093 allmänhet 42
6094 allmänheten 47
6095 allmänhetens 15
6096 allmänintresse 1
6097 allmänna 132
6098 allmännas 1
6099 allmänne 1
6100 allmännyttig 2
6101 allmännyttiga 7
6102 allmänpolitisk 1
6103 allmänt 56
6104 allokeringar 1
6105 allomfattande 1
6106 allra 40
6107 alls 75
6108 allsidig 2
6109 allsidigt 2
6110 allsmäktighet 1
6111 allt 617
6112 allteftersom 7
6113 alltfler 3
6114 alltför 133
6115 alltid 210
6116 alltifrån 3
6117 alltihop 15
6118 allting 18
6119 alltjämt 7
6120 alltmer 13
6121 alltsammans 10
6122 alltsedan 4
6123 alltså 191
6124 allvar 36
6125 allvaret 3
6126 allvarlig 37
6127 allvarliga 80
6128 allvarligare 11
6129 allvarligaste 6
6130 allvarligt 64
6131 allvarsamt 1
6132 alster 1
6133 alt 1
6134 altare 1
6135 alternativ 28
6136 alternativa 7
6137 alternativen 1
6138 alternativet 3
6139 alternativt 1
6140 amatördiplomati 1
6141 ambassad 1
6142 ambassadör 2
6143 ambassadören 1
6144 ambassadörer 3
6145 ambition 17
6146 ambitionen 7
6147 ambitioner 25
6148 ambitionerna 1
6149 ambitionernas 2
6150 ambitiös 18
6151 ambitiösa 22
6152 ambitiösare 2
6153 ambitiöse 1
6154 ambitiöst 10
6155 ambulans 1
6156 ambulanser 1
6157 amerikan 1
6158 amerikanarna 1
6159 amerikanen 1
6160 amerikaner 1
6161 amerikanerna 14
6162 amerikansk 5
6163 amerikanska 51
6164 amerikanske 1
6165 amerikanskt 2
6166 amfiteatraliskt 1
6167 amiraler 1
6168 ammunition 1
6169 an 20
6170 ana 7
6171 anade 2
6172 analogt 1
6173 analys 40
6174 analysen 10
6175 analyser 4
6176 analysera 21
6177 analyserar 1
6178 analyseras 5
6179 analyserat 3
6180 analyserna 1
6181 analytiskt 2
6182 anamma 3
6183 anammande 1
6184 anammar 1
6185 anammat 4
6186 anammats 1
6187 anar 1
6188 anblick 1
6189 anblicken 3
6190 anbudsförfarande 1
6191 anbudsförfaranden 1
6192 anbudsförfarandet 2
6193 anbudsgivare 1
6194 anbudsgivningen 1
6195 anbudsinfordran 2
6196 and 9
6197 anda 23
6198 andades 2
6199 andaluser 2
6200 andalusier 3
6201 andalusierna 1
6202 andalusiska 1
6203 andan 10
6204 andas 3
6205 ande 1
6206 andedräkt 1
6207 andel 15
6208 andelar 4
6209 andelen 7
6210 andemening 2
6211 andemeningen 5
6212 andens 1
6213 andetag 2
6214 andfådd 1
6215 andhämtningens 1
6216 andlig 1
6217 andliga 3
6218 andlige 1
6219 andra 1089
6220 andrabehandling 1
6221 andrabehandlingsrekommendation 5
6222 andrabehandlingsrekommendationen 5
6223 andrahandsbehandlingsrekommendation 1
6224 andrakammare 1
6225 andras 7
6226 andre 4
6227 andres 1
6228 anemi 1
6229 anfall 2
6230 anfallen 2
6231 anföra 4
6232 anförande 21
6233 anföranden 15
6234 anförandena 3
6235 anförandet 3
6236 anföras 1
6237 anförs 2
6238 anfört 2
6239 anförtro 1
6240 anförtros 3
6241 anförtrott 1
6242 anförtrotts 2
6243 angav 3
6244 angavs 2
6245 ange 19
6246 angelägen 14
6247 angelägenhet 11
6248 angelägenheten 3
6249 angelägenheter 11
6250 angelägenheterna 1
6251 angeläget 9
6252 angelägna 12
6253 angelägnare 1
6254 angenäm 3
6255 angenämt 1
6256 anger 17
6257 anges 31
6258 angetts 2
6259 angivandet 2
6260 angivare 2
6261 angivarna 1
6262 angivelse 1
6263 angiven 1
6264 angiveri 1
6265 angivit 4
6266 angivna 2
6267 angjorde 1
6268 anglosaxiska 1
6269 angolaner 1
6270 angolanska 10
6271 angrep 2
6272 angrepp 9
6273 angreppen 1
6274 angreppet 1
6275 angreppskrig 1
6276 angreppssätt 4
6277 angripa 13
6278 angripas 2
6279 angripen 2
6280 angriper 4
6281 angrips 1
6282 angränsande 5
6283 angående 72
6284 angår 6
6285 angör 1
6286 anhängare 8
6287 anhängiggjort 1
6288 anhängiggöranden 1
6289 anhålla 2
6290 anhållnas 1
6291 anhållne 1
6292 anhöriga 2
6293 aning 12
6294 aningar 1
6295 aningen 2
6296 aningslösa 1
6297 ankar 3
6298 ankare 1
6299 ankaret 2
6300 ankarplats 1
6301 anklaga 1
6302 anklagad 1
6303 anklagade 4
6304 anklagades 2
6305 anklagas 4
6306 anklagelse 1
6307 anklagelsen 1
6308 anklagelser 6
6309 anklagelserna 6
6310 anklarna 1
6311 anknutna 1
6312 anknytning 4
6313 anknyts 1
6314 ankommer 1
6315 ankomst 2
6316 ankomsten 1
6317 ankrade 2
6318 anlag 1
6319 anlagd 2
6320 anlagda 1
6321 anlagt 2
6322 anlagts 1
6323 anledning 77
6324 anledningar 9
6325 anledningarna 2
6326 anledningen 52
6327 anletsdrag 1
6328 anlitat 1
6329 anlägga 1
6330 anlägger 2
6331 anläggning 6
6332 anläggningar 5
6333 anläggningarna 2
6334 anläggningarnas 1
6335 anläggningen 3
6336 anläggningsarbeten 1
6337 anläggs 1
6338 anlända 2
6339 anlände 2
6340 anländer 1
6341 anlänt 2
6342 anlöpa 1
6343 anlöper 5
6344 anmodade 3
6345 anmodan 1
6346 anmodar 1
6347 anmäla 4
6348 anmälan 4
6349 anmälda 2
6350 anmäler 1
6351 anmälning 1
6352 anmälningar 2
6353 anmälningsplikt 3
6354 anmälningsplikten 1
6355 anmälningsplikter 1
6356 anmälningssystemet 3
6357 anmäls 2
6358 anmält 3
6359 anmälts 1
6360 anmärkning 13
6361 anmärkningar 8
6362 anmärkningarna 2
6363 anmärkningen 1
6364 anmärkningsvärd 2
6365 anmärkningsvärda 4
6366 anmärkningsvärt 6
6367 annalkande 2
6368 annan 154
6369 annanstans 6
6370 annars 30
6371 annat 269
6372 annonsera 1
6373 annorlunda 23
6374 annorstädes 4
6375 anomali 1
6376 anonym 2
6377 anonyma 2
6378 anonymitet 1
6379 anordna 3
6380 anordnade 5
6381 anordnas 2
6382 anordnats 1
6383 anordning 4
6384 anordningar 3
6385 anpassa 25
6386 anpassad 9
6387 anpassade 9
6388 anpassas 14
6389 anpassat 5
6390 anpassats 1
6391 anpassbarhet 1
6392 anpassning 14
6393 anpassningar 5
6394 anpassningarna 3
6395 anpassningen 6
6396 anpassningsbarhet 2
6397 anpassningsetappen 1
6398 anpassningsfasen 1
6399 anpassningsförmåga 4
6400 anpassningsproblem 1
6401 anropa 1
6402 anrätta 1
6403 ansade 1
6404 ansamlingen 1
6405 ansats 4
6406 ansatsen 2
6407 ansatser 5
6408 ansatserna 1
6409 anse 10
6410 ansedda 1
6411 anseende 9
6412 ansenlig 3
6413 ansenliga 1
6414 ansenligt 1
6415 anser 494
6416 anses 24
6417 ansett 7
6418 ansikte 27
6419 ansikten 6
6420 ansiktena 3
6421 ansiktet 10
6422 ansiktshuden 1
6423 ansiktslöse 1
6424 ansiktsuttryck 1
6425 ansjovis 4
6426 ansjovisbestånden 6
6427 ansjovisbeståndet 3
6428 ansjovisen 1
6429 ansjovisfiske 1
6430 ansjovisfisket 2
6431 ansjoviskvoten 1
6432 ansjoviskvoter 1
6433 anskaffat 1
6434 anskaffning 2
6435 anskrämliga 1
6436 anslag 26
6437 anslagen 20
6438 anslaget 6
6439 anslagits 1
6440 anslagna 2
6441 anslagsbeviljandet 1
6442 anslagsförbrukning 1
6443 anslagsfördelningen 1
6444 anslogs 1
6445 ansluta 30
6446 anslutande 1
6447 anslutas 1
6448 ansluter 17
6449 anslutit 5
6450 anslutits 1
6451 anslutna 3
6452 anslutning 39
6453 anslutningar 1
6454 anslutningen 18
6455 anslutningsfil 18
6456 anslutningsfilen 9
6457 anslutningsfilens 1
6458 anslutningsfiler 1
6459 anslutningsförfarandet 3
6460 anslutningsförhandlingarna 6
6461 anslutningsinformationen 5
6462 anslutningsländerna 1
6463 anslutningsmedel 1
6464 anslutningsprocess 1
6465 anslutningsprojektet 1
6466 anslutningsstrategin 1
6467 ansluts 2
6468 anslå 4
6469 anslår 2
6470 anslås 4
6471 anslöt 2
6472 anspelade 2
6473 anspelningar 1
6474 anspråk 14
6475 anspråksfulla 1
6476 anspråkslösa 2
6477 anspråkslösaste 1
6478 anspråkslöshet 1
6479 anstrykning 1
6480 anstränga 8
6481 ansträngda 1
6482 ansträngde 4
6483 anstränger 10
6484 ansträngning 8
6485 ansträngningar 75
6486 ansträngningarna 11
6487 ansträngs 1
6488 ansträngt 5
6489 anställa 8
6490 anställande 1
6491 anställbara 1
6492 anställbarhet 6
6493 anställbarheten 2
6494 anställd 3
6495 anställda 38
6496 anställdas 8
6497 anställer 1
6498 anställning 10
6499 anställningarna 2
6500 anställningsförhållanden 1
6501 anställningskontrakt 1
6502 anställningsmöjligheter 1
6503 anställningsvillkor 1
6504 anställt 1
6505 anställts 1
6506 anständig 4
6507 anständiga 5
6508 anständighet 3
6509 anständigt 3
6510 anstår 1
6511 ansvar 219
6512 ansvara 6
6513 ansvarar 13
6514 ansvaret 76
6515 ansvarig 38
6516 ansvariga 52
6517 ansvarige 3
6518 ansvarigt 6
6519 ansvarsavgränsning 1
6520 ansvarsbefrielse 1
6521 ansvarsbefrielsen 1
6522 ansvarsbördor 1
6523 ansvarsfrihet 34
6524 ansvarsfriheten 7
6525 ansvarsfrihetsrapport 1
6526 ansvarsfrågan 3
6527 ansvarsfrågorna 1
6528 ansvarsfull 3
6529 ansvarsfulla 6
6530 ansvarsfullt 11
6531 ansvarsfyllda 1
6532 ansvarsfördelning 2
6533 ansvarsfördelningen 3
6534 ansvarsförhållandena 1
6535 ansvarskultur 1
6536 ansvarskännande 2
6537 ansvarskänsla 3
6538 ansvarsområde 7
6539 ansvarsområden 3
6540 ansvarsområdena 1
6541 ansvarsområdet 1
6542 ansvarsordning 1
6543 ansvarsposter 4
6544 ansvarstagande 2
6545 ansvarstagandet 1
6546 ansvarstilldelning 1
6547 ansvarsuppgifter 1
6548 ansåg 18
6549 ansågs 5
6550 ansöka 2
6551 ansökan 12
6552 ansökande 2
6553 ansökarland 2
6554 ansökarländer 4
6555 ansökarländerna 12
6556 ansöker 2
6557 ansökningar 3
6558 ansökningsbestämmelser 1
6559 ansökt 2
6560 anta 58
6561 antagande 8
6562 antaganden 2
6563 antagandeprocessen 1
6564 antagandet 20
6565 antagen 3
6566 antagit 25
6567 antagits 20
6568 antagligen 10
6569 antagna 6
6570 antal 139
6571 antalet 66
6572 antar 23
6573 antas 26
6574 ante 5
6575 ante-systemet 1
6576 antecknade 2
6577 antecknat 1
6578 anteckningsblock 1
6579 anteckningsbok 2
6580 anteckningsboken 1
6581 antenner 2
6582 anti-europeisk 1
6583 anti-europeiska 1
6584 anti-gemenskapliga 1
6585 anti-irländska 1
6586 anti-rasistiska 1
6587 antibedrägerilagstiftning 1
6588 antibiotika 7
6589 antibiotikaresistensens 1
6590 antibiotikum 1
6591 antidemokratiska 1
6592 antidiskrimineringslagar 1
6593 antieuropeiska 2
6594 antifascist 1
6595 antifascistiska 2
6596 antifolklig 1
6597 antika 2
6598 antikaffär 1
6599 antikens 1
6600 antikolonialism 1
6601 antikryptogam 2
6602 antimögelmedel 1
6603 antingen 25
6604 antipersonella 2
6605 antisemitiska 1
6606 antisemitism 3
6607 antisociala 1
6608 antiterroristoperation 1
6609 antites 1
6610 antitrustbestämmelserna 1
6611 antog 42
6612 antogs 22
6613 antropogenisk 1
6614 antropolog 1
6615 antyda 2
6616 antydan 3
6617 antydas 1
6618 antydde 4
6619 antyddes 1
6620 antyder 6
6621 antytt 1
6622 antågande 1
6623 anvisade 1
6624 anvisning 1
6625 anvisningar 2
6626 anvisningarna 2
6627 använd 3
6628 använda 135
6629 användande 4
6630 användandet 1
6631 användare 9
6632 användaren 3
6633 användarens 1
6634 användares 2
6635 användargränssnitt 1
6636 användargränssnittet 3
6637 användarkrav 1
6638 användarkraven 1
6639 användarna 4
6640 användarnas 3
6641 användas 66
6642 användbar 4
6643 användbara 4
6644 användbarhet 1
6645 användbart 7
6646 använde 14
6647 använder 68
6648 användes 7
6649 användning 44
6650 användningarna 1
6651 användningen 33
6652 används 62
6653 använt 12
6654 använts 13
6655 apartheid 1
6656 apartheid-ordning 1
6657 apos 1
6658 apostrof 1
6659 apotek 1
6660 apoteket 1
6661 apparat 1
6662 apparaten 1
6663 apparater 2
6664 apparaterna 1
6665 appell 1
6666 appellationsdomstolen 1
6667 applåder 15
6668 applådera 1
6669 applåderade 1
6670 applåderar 3
6671 april 21
6672 apropå 3
6673 aptit 1
6674 arab 1
6675 arabisk 1
6676 arabisk-israeliska 1
6677 arabiska 11
6678 arabstat 1
6679 arabstater 1
6680 arabvärlden 1
6681 arbeta 117
6682 arbetad 1
6683 arbetade 10
6684 arbetande 5
6685 arbetar 68
6686 arbetare 10
6687 arbetaren 1
6688 arbetarens 1
6689 arbetarklassens 1
6690 arbetarna 3
6691 arbetarnas 2
6692 arbetarpartis 1
6693 arbetarstadsdelar 1
6694 arbetas 1
6695 arbetat 30
6696 arbete 272
6697 arbeten 17
6698 arbetena 2
6699 arbetet 81
6700 arbetets 2
6701 arbets- 3
6702 arbetsanda 1
6703 arbetsaspekter 1
6704 arbetsavtal 2
6705 arbetsbelastning 1
6706 arbetsbeskrivningar 1
6707 arbetsbörda 4
6708 arbetsbördan 1
6709 arbetsdokument 4
6710 arbetsdokumenten 1
6711 arbetsformer 2
6712 arbetsfrågorna 1
6713 arbetsfördelning 2
6714 arbetsförhållanden 2
6715 arbetsförmedlingar 1
6716 arbetsförmedlingen 1
6717 arbetsförmåga 1
6718 arbetsgivare 10
6719 arbetsgivaren 2
6720 arbetsgivarens 2
6721 arbetsgivarna 2
6722 arbetsgivarnas 3
6723 arbetsgivarorganisationen 1
6724 arbetsgivarparti 1
6725 arbetsgrupp 17
6726 arbetsgruppen 3
6727 arbetsgrupper 4
6728 arbetsinkomster 1
6729 arbetsinsats 3
6730 arbetsinsatser 2
6731 arbetsinsatserna 1
6732 arbetsintensiva 2
6733 arbetskontraktet 1
6734 arbetskraft 14
6735 arbetskraften 7
6736 arbetskraftens 1
6737 arbetskraftsintensiva 2
6738 arbetskraftsrörlighet 1
6739 arbetskultur 2
6740 arbetskvalitet 2
6741 arbetslagstiftning 1
6742 arbetsliv 4
6743 arbetslivet 9
6744 arbetslivets 1
6745 arbetslösa 21
6746 arbetslösas 2
6747 arbetslöshet 36
6748 arbetslösheten 66
6749 arbetslöshetens 3
6750 arbetslöshetsersättningen 1
6751 arbetslöshetsnivåer 1
6752 arbetslöshetspolitik 1
6753 arbetslöshetsproblemet 2
6754 arbetslöshetssiffrorna 3
6755 arbetslöshetsunderstöd 1
6756 arbetsmarknad 8
6757 arbetsmarknaden 38
6758 arbetsmarknadens 16
6759 arbetsmarknaderna 2
6760 arbetsmarknadsfrågor 1
6761 arbetsmarknadsförhållandena 1
6762 arbetsmarknadslagarna 1
6763 arbetsmarknadsministern 1
6764 arbetsmarknadsministrar 1
6765 arbetsmarknadsmyndigheter 1
6766 arbetsmarknadsorganisationerna 1
6767 arbetsmarknadsparternas 1
6768 arbetsmarknadspolitik 1
6769 arbetsmarknadspolitiken 4
6770 arbetsmarknadsproblem 1
6771 arbetsmetod 2
6772 arbetsmetoden 2
6773 arbetsmetoder 4
6774 arbetsmetoderna 3
6775 arbetsmigration 1
6776 arbetsmiljö 1
6777 arbetsmotivation 1
6778 arbetsmängd 1
6779 arbetsmässiga 1
6780 arbetsmöjligheter 1
6781 arbetsnormer 3
6782 arbetsnormerna 1
6783 arbetsoduglig 1
6784 arbetsområdet 2
6785 arbetsordning 4
6786 arbetsordningen 22
6787 arbetsorganisation 2
6788 arbetsorganisationen 2
6789 arbetsorganiseringen 1
6790 arbetsperiod 1
6791 arbetsplan 1
6792 arbetsplanen 5
6793 arbetsplaner 1
6794 arbetsplats 1
6795 arbetsplatsen 3
6796 arbetsplatser 14
6797 arbetsplatserna 2
6798 arbetsplikt 1
6799 arbetspost 1
6800 arbetsprocessen 1
6801 arbetsprogram 13
6802 arbetsprogrammet 4
6803 arbetsrelationerna 1
6804 arbetsrum 1
6805 arbetsrutiner 1
6806 arbetsrätt 1
6807 arbetsrätten 1
6808 arbetsrättsliga 1
6809 arbetssammanträde 1
6810 arbetsskapande 1
6811 arbetsstyrka 2
6812 arbetsstyrkan 1
6813 arbetssystem 1
6814 arbetssätt 1
6815 arbetssättet 1
6816 arbetssökande 1
6817 arbetstagare 46
6818 arbetstagaren 5
6819 arbetstagarens 1
6820 arbetstagares 4
6821 arbetstagarna 22
6822 arbetstagarnas 11
6823 arbetstid 2
6824 arbetstiden 6
6825 arbetstidens 1
6826 arbetstider 2
6827 arbetstidsdirektivet 2
6828 arbetstidsförkortning 3
6829 arbetstidskriterierna 1
6830 arbetstidsordning 1
6831 arbetstidsreglerna 1
6832 arbetstidsutformning 1
6833 arbetstillfällen 94
6834 arbetstillfällena 4
6835 arbetstillstånd 5
6836 arbetstillståndet 1
6837 arbetsuppgifter 4
6838 arbetsverktyg 1
6839 arbetsvillkor 7
6840 arbetsvillkoren 4
6841 arbetsvärlden 1
6842 arbetsyta 2
6843 are 1
6844 arena 1
6845 arenan 1
6846 argent 1
6847 argument 28
6848 argumentation 1
6849 argumentationen 1
6850 argumentationskraft 1
6851 argumenten 5
6852 argumentera 3
6853 argumenterar 3
6854 argumentet 4
6855 aristokrat 1
6856 arkeolog 1
6857 arkeologiska 1
6858 arkitekter 1
6859 arkitektur 1
6860 arkiv 1
6861 arkiveras 1
6862 arkivutrymmen 1
6863 arm 3
6864 armar 4
6865 armarna 2
6866 armarnas 1
6867 armbandsur 1
6868 armbågarna 1
6869 armbåge 1
6870 armbågen 1
6871 armen 2
6872 armenierna 2
6873 armod 2
6874 armé 8
6875 armén 4
6876 arméns 2
6877 arrangemang 6
6878 arrangemangen 2
6879 arrangera 3
6880 arrangerandet 1
6881 arrangerat 1
6882 arrest 1
6883 arresterad 2
6884 arresterades 6
6885 arresterats 1
6886 arresteringar 3
6887 arrogans 1
6888 arrogant 1
6889 arroganta 2
6890 arsenal 1
6891 art 13
6892 arte 1
6893 artefakt 1
6894 arten 2
6895 arter 9
6896 arterna 3
6897 artificiell 1
6898 artificiella 1
6899 artig 1
6900 artiga 2
6901 artighet 3
6902 artighetsgest 1
6903 artikel 234
6904 artikeln 1
6905 artiklar 10
6906 artiklarna 11
6907 artister 1
6908 arton 5
6909 artonhundratalet 1
6910 artonhundratalsstil 1
6911 artärer 1
6912 arv 13
6913 arven 1
6914 arvet 3
6915 arvode 1
6916 arvoden 1
6917 arvsynden 1
6918 as 1
6919 asfalterade 1
6920 asiatiska 1
6921 ask 1
6922 aska 2
6923 askar 1
6924 asken 1
6925 askenasernas 1
6926 asket 1
6927 askkoppar 1
6928 asocial 1
6929 aspekt 18
6930 aspekten 15
6931 aspekter 51
6932 aspekterna 10
6933 aspirera 1
6934 assegajer 1
6935 assimilering 1
6936 assistans 1
6937 assistent 2
6938 assistenter 2
6939 assistenterna 4
6940 assistentstadga 1
6941 assisterad 1
6942 assistito 1
6943 associerade 4
6944 associeras 1
6945 associering 1
6946 associeringsavtal 9
6947 associeringsavtalen 2
6948 associeringsavtalet 6
6949 associeringsförfarande 1
6950 associeringsprocessen 2
6951 asterisk 1
6952 asteroid 1
6953 asteroiden 1
6954 astma 1
6955 astronomen 1
6956 astronomiska 1
6957 asyl 10
6958 asyl- 2
6959 asylbeslut 1
6960 asylfrågan 1
6961 asylförfarande 2
6962 asylförfarandet 1
6963 asylpolitik 1
6964 asylrätt 4
6965 asylsökande 18
6966 asylsökandena 1
6967 asymmetrierna 1
6968 asymmetriska 1
6969 at 2
6970 ateister 1
6971 atlantalliansen 1
6972 atlantfart 1
6973 atlantkusten 1
6974 atmosfär 5
6975 atmosfärens 1
6976 atomenergimyndigheten 1
6977 atomenergiorganet 2
6978 atomforskningscentret 1
6979 atomkraften 1
6980 att 18791
6981 attack 2
6982 attacken 1
6983 attacker 7
6984 attackerna 1
6985 attentat 3
6986 attentatet 1
6987 attesterats 1
6988 attityd 15
6989 attityder 2
6990 attraktionskraft 1
6991 attraktiv 2
6992 attraktiva 3
6993 attraktivt 2
6994 attributen 1
6995 atypiska 1
6996 atypiskt 1
6997 auctoritas 1
6998 audio-visuella 1
6999 audiovisuella 1
7000 auditorium 1
7001 augusti 5
7002 auktionerna 1
7003 auktorisation 3
7004 auktoriserad 1
7005 auktoriserade 1
7006 auktoriseringar 1
7007 auktoritativ 1
7008 auktoritet 7
7009 auktoriteter 1
7010 automatik 2
7011 automatisk 1
7012 automatiska 2
7013 automatiskt 20
7014 autonoma 2
7015 autonomi 3
7016 autonomin 1
7017 autopilot 1
7018 av 8457
7019 avancera 2
7020 avancerade 1
7021 avancerat 2
7022 avant 2
7023 avart 1
7024 avbetalning 1
7025 avbrott 4
7026 avbrottet 5
7027 avbruten 3
7028 avbrutits 2
7029 avbrutna 1
7030 avbryta 2
7031 avbryter 5
7032 avbryts 2
7033 avbröt 11
7034 avbröts 13
7035 avböjer 1
7036 avdela 4
7037 avdelar 1
7038 avdelning 11
7039 avdelningar 4
7040 avdelningarna 1
7041 avdelningen 2
7042 avdelnings- 1
7043 avdemokratiserar 1
7044 avec 2
7045 avenyn 1
7046 aversion 1
7047 aveuropeisering 1
7048 avfall 39
7049 avfallet 15
7050 avfallets 1
7051 avfalls- 1
7052 avfallsdirektiven 1
7053 avfallsfisk 1
7054 avfallshantering 2
7055 avfallshanteringen 2
7056 avfallshanteringens 1
7057 avfallshanteringsavgift 1
7058 avfallsinsamlaren 1
7059 avfallsmängd 1
7060 avfallsström 1
7061 avfallsströmmar 2
7062 avfallsströmmarna 1
7063 avfallssystem 1
7064 avfallsämnen 1
7065 avfolkas 1
7066 avfolkats 1
7067 avfolkning 3
7068 avfolkningsbygder 1
7069 avfolkningsvåg 1
7070 avfälliga 1
7071 avfärd 1
7072 avfärdad 1
7073 avfärdade 2
7074 avförd 1
7075 avfördes 1
7076 avförs 1
7077 avförts 1
7078 avgaser 1
7079 avgav 2
7080 avge 6
7081 avger 6
7082 avges 1
7083 avgett 1
7084 avgick 4
7085 avgift 4
7086 avgifter 8
7087 avgiftsutjämning 1
7088 avgivit 1
7089 avgivits 1
7090 avgjorde 2
7091 avgjort 3
7092 avgjorts 2
7093 avgrund 1
7094 avgränsa 1
7095 avgränsade 3
7096 avgränsar 1
7097 avgränsat 1
7098 avgå 2
7099 avgående 1
7100 avgång 6
7101 avgångsåtgärder 1
7102 avgår 1
7103 avgått 1
7104 avgör 5
7105 avgöra 19
7106 avgörande 113
7107 avgörandet 2
7108 avgöras 4
7109 avgörs 5
7110 avhandla 1
7111 avhandlas 2
7112 avhandlats 1
7113 avhjälpa 3
7114 avhjälpande 1
7115 avhjälpas 1
7116 avhjälps 1
7117 avhjälpts 2
7118 avhänder 1
7119 avhängig 2
7120 avhängigt 2
7121 avhålla 2
7122 avhållit 1
7123 avigsidor 1
7124 aviserade 3
7125 aviserar 2
7126 aviseras 1
7127 aviserat 2
7128 aviserats 2
7129 avisering 1
7130 avkall 2
7131 avkastning 5
7132 avkastningen 3
7133 avkastningsdjur 1
7134 avklarad 2
7135 avklarats 1
7136 avkrok 1
7137 avkrävas 2
7138 avkrävt 1
7139 avkunnar 2
7140 avlade 2
7141 avlagd 1
7142 avlagt 1
7143 avlastning 1
7144 avledda 2
7145 avleder 1
7146 avlida 1
7147 avlivad 1
7148 avlivar 1
7149 avlivas 1
7150 avlivning 1
7151 avloppet 2
7152 avloppshål 1
7153 avloppsrör 1
7154 avlutat 1
7155 avlyssna 1
7156 avlyssnas 1
7157 avlyssning 11
7158 avlyssningen 4
7159 avlyssningssystemet 1
7160 avlägga 2
7161 avlägsen 5
7162 avlägset 6
7163 avlägsna 22
7164 avlägsnade 2
7165 avlägsnande 2
7166 avlägsnandet 2
7167 avlägsnas 1
7168 avlägsnat 1
7169 avlämnats 1
7170 avlöses 1
7171 avlösning 1
7172 avmagringskur 1
7173 avmattning 2
7174 avnjöt 1
7175 avocadokärnan 1
7176 avocat 2
7177 avoghet 1
7178 avogt 1
7179 avpassade 1
7180 avprickning 1
7181 avrapportering 1
7182 avreglera 4
7183 avreglerad 5
7184 avreglerade 2
7185 avreglerar 2
7186 avregleras 2
7187 avreglerat 2
7188 avreglering 39
7189 avregleringar 1
7190 avregleringen 44
7191 avregleringens 1
7192 avregleringsetapp 3
7193 avregleringsfas 1
7194 avregleringsområdet 1
7195 avregleringspolitiken 1
7196 avregleringsprocess 1
7197 avregleringsprocessen 1
7198 avregleringsscenarierna 1
7199 avregleringssteget 1
7200 avresan 1
7201 avrinningsområde 1
7202 avrinningsområden 1
7203 avrunda 1
7204 avrätta 1
7205 avrättades 1
7206 avrättat 1
7207 avråda 1
7208 avröjda 1
7209 avsaknad 5
7210 avsaknaden 14
7211 avsatsen 2
7212 avsatt 3
7213 avsatta 3
7214 avsattes 2
7215 avsatts 3
7216 avse 4
7217 avsedd 9
7218 avsedda 13
7219 avseende 70
7220 avseenden 19
7221 avseendena 1
7222 avseendet 42
7223 avser 63
7224 avses 9
7225 avsett 16
7226 avsevärd 6
7227 avsevärda 11
7228 avsevärt 15
7229 avsides 3
7230 avsikt 62
7231 avsikten 11
7232 avsikter 16
7233 avsikterna 3
7234 avsiktlig 2
7235 avsiktliga 3
7236 avsiktligt 4
7237 avsiktsförklaring 1
7238 avsiktsförklaringar 2
7239 avskaffa 23
7240 avskaffade 3
7241 avskaffades 2
7242 avskaffande 4
7243 avskaffandet 3
7244 avskaffar 4
7245 avskaffas 1
7246 avskaffat 1
7247 avskaffats 1
7248 avsked 2
7249 avskeda 2
7250 avskedande 1
7251 avskedar 1
7252 avskedat 1
7253 avskilda 1
7254 avskiljas 1
7255 avskriva 1
7256 avskrivning 1
7257 avskruvad 1
7258 avskräcka 3
7259 avskräckande 2
7260 avskräckning 1
7261 avskräcks 1
7262 avskrädeshög 1
7263 avskuren 1
7264 avsky 4
7265 avskydd 1
7266 avskydde 1
7267 avskyr 1
7268 avskytt 1
7269 avskyvärda 3
7270 avskyvärt 1
7271 avskärma 2
7272 avskärmar 1
7273 avskärmat 1
7274 avskärmning 1
7275 avslag 2
7276 avslitet 1
7277 avslog 6
7278 avslogs 3
7279 avsluta 37
7280 avslutad 68
7281 avslutade 11
7282 avslutades 12
7283 avslutande 5
7284 avslutandet 1
7285 avslutar 10
7286 avslutas 12
7287 avslutat 9
7288 avslutats 4
7289 avslutning 6
7290 avslutningen 2
7291 avslutningsvis 13
7292 avslängd 1
7293 avslå 3
7294 avslår 1
7295 avslås 2
7296 avslöja 2
7297 avslöjade 3
7298 avslöjades 1
7299 avslöjande 3
7300 avslöjanden 1
7301 avslöjar 9
7302 avslöjas 1
7303 avslöjat 1
7304 avsmak 3
7305 avsmalnande 1
7306 avsnitt 7
7307 avsnitten 2
7308 avsnittet 4
7309 avspegla 1
7310 avspeglar 6
7311 avspeglas 7
7312 avspänd 1
7313 avspända 1
7314 avspänning 1
7315 avspärrningar 1
7316 avstamp 1
7317 avstannat 1
7318 avsteg 1
7319 avstod 6
7320 avstänga 1
7321 avstängde 1
7322 avstängning 2
7323 avstå 16
7324 avståenden 1
7325 avstånd 16
7326 avstånden 2
7327 avståndet 10
7328 avståndstagande 3
7329 avstår 7
7330 avstått 8
7331 avsägande 1
7332 avsätta 6
7333 avsättas 1
7334 avsätter 1
7335 avsättningarna 1
7336 avsåg 6
7337 avtacklade 1
7338 avtal 126
7339 avtalade 3
7340 avtalas 1
7341 avtalat 3
7342 avtalats 4
7343 avtalen 22
7344 avtalens 1
7345 avtalet 70
7346 avtalets 7
7347 avtals 1
7348 avtalsförbindelser 1
7349 avtalsinnehållet 1
7350 avtalslösning 1
7351 avtalspart 1
7352 avtalsparterna 2
7353 avtalsslutande 1
7354 avtalstexten 1
7355 avtalstexterna 1
7356 avtalsvillkoren 2
7357 avtar 1
7358 avtecknade 4
7359 avtecknat 1
7360 avtvinga 1
7361 avund 1
7362 avundades 1
7363 avundas 2
7364 avundsjuka 1
7365 avundsvärda 1
7366 avvakta 5
7367 avvaktan 6
7368 avvaktande 2
7369 avvaktar 3
7370 avveckla 6
7371 avvecklas 4
7372 avvecklat 2
7373 avvecklats 1
7374 avveckling 3
7375 avverkningsklara 1
7376 avvika 1
7377 avvikande 4
7378 avvikelse 1
7379 avvikelser 4
7380 avviker 3
7381 avvisa 9
7382 avvisade 3
7383 avvisades 1
7384 avvisande 1
7385 avvisandet 1
7386 avvisar 6
7387 avvisas 1
7388 avvisat 3
7389 avvisats 2
7390 avvisning 2
7391 avvägd 4
7392 avvägning 4
7393 avvägningar 1
7394 avvägningen 1
7395 avvägningsfall 1
7396 avvägs 1
7397 avvägt 1
7398 avväpnade 1
7399 avvärja 3
7400 avyttring 1
7401 axeln 3
7402 axelryckning 3
7403 axla 1
7404 axlar 3
7405 axlarna 6
7406 b 8
7407 baby 1
7408 babyn 1
7409 bacill 1
7410 back-position 1
7411 backa 1
7412 backade 4
7413 backen 2
7414 backshish-mentalitet 1
7415 bad 15
7416 bada 1
7417 badar 1
7418 badet 1
7419 badhytterna 1
7420 badkaret 1
7421 badrummet 3
7422 badwill 1
7423 bagage 1
7424 bagaget 1
7425 bagatell 1
7426 bagatelliserar 1
7427 bagatellisering 1
7428 bain 1
7429 bak 5
7430 bakat 1
7431 bakbundna 1
7432 bakdanta 1
7433 bakdörren 4
7434 baken 1
7435 bakficka 1
7436 bakfönstret 1
7437 bakgata 1
7438 bakgrund 70
7439 bakgrunden 14
7440 bakgrundsförslag 1
7441 bakgrundsnivå 1
7442 bakgrundsutsläpp 1
7443 bakgrundsvärdena 2
7444 bakgård 1
7445 bakgårdar 1
7446 bakhåll 1
7447 bakifrån 2
7448 bakning 1
7449 bakom 95
7450 bakomliggande 6
7451 bakre 1
7452 baksidestext 1
7453 bakslag 1
7454 bakslaget 1
7455 bakslugt 1
7456 baksätet 3
7457 baktalade 1
7458 baktanken 1
7459 bakvägen 1
7460 bakvägspolitik 1
7461 bakåt 6
7462 bakåtsträvande 2
7463 bakåtverkande 1
7464 balans 45
7465 balansen 14
7466 balanser 2
7467 balansera 3
7468 balanserad 15
7469 balanserade 6
7470 balanserande 1
7471 balanserar 2
7472 balanseras 1
7473 balanserat 8
7474 balansering 1
7475 balansräkningar 1
7476 balansövning 1
7477 baldakinförsedda 1
7478 balen 3
7479 balkan 1
7480 ballader 1
7481 ballast 1
7482 ballon 1
7483 baltiska 1
7484 bana 4
7485 banalisera 2
7486 banaliserar 1
7487 banaliseringen 1
7488 bananerna 1
7489 bananrepubliker 1
7490 banar 1
7491 banat 1
7492 banbrytande 1
7493 band 17
7494 banden 3
7495 banderoll 2
7496 bandet 2
7497 banditer 1
7498 bank 3
7499 banka 1
7500 bankade 1
7501 banken 1
7502 bankens 1
7503 banker 4
7504 banketter 1
7505 bankförvaltningen 1
7506 bankgarantier 5
7507 bankirer 2
7508 bankkoncernerna 1
7509 bankkonton 2
7510 bankrutt 2
7511 banksekretessen 1
7512 banksystemet 1
7513 bannlysningen 1
7514 bannlysts 1
7515 banor 3
7516 bantas 1
7517 bantning 1
7518 bantningen 1
7519 bantningskur 1
7520 bar 16
7521 bara 861
7522 baracker 1
7523 barbari 1
7524 barbariet 2
7525 barbariets 1
7526 barbariska 2
7527 barbariskt 1
7528 barberarna 1
7529 baren 2
7530 barens 1
7531 barerna 1
7532 barkborren 1
7533 barm 2
7534 barn 64
7535 barn- 1
7536 barnadödlighet 4
7537 barnadödligheten 1
7538 barnafödande 1
7539 barnbarn 1
7540 barnbedrägeri 1
7541 barndom 1
7542 barndomen 1
7543 barndödlighet 3
7544 barndödligheten 1
7545 barnen 10
7546 barnens 8
7547 barnet 3
7548 barnets 1
7549 barnhandel 1
7550 barnhälsoproblemet 1
7551 barnmorska 1
7552 barnomsorg 2
7553 barnpornografi 2
7554 barns 5
7555 barnsligaste 1
7556 barnungar 1
7557 baron 1
7558 barriärer 2
7559 bars 2
7560 barskt 1
7561 bart 1
7562 bartender 1
7563 bas 6
7564 basackompanjemanget 1
7565 basar 2
7566 base 1
7567 baseball 1
7568 baseballmössor 1
7569 baseballresultaten 1
7570 basen 4
7571 baser 1
7572 basera 2
7573 baserad 5
7574 baserade 6
7575 baserar 4
7576 baseras 14
7577 baserat 4
7578 basförsörjning 1
7579 basis 6
7580 bask 4
7581 baskisk 3
7582 baskiska 12
7583 baskiskt 1
7584 baskolumnens 1
7585 baskrar 1
7586 basnivå 1
7587 bastardhunden 1
7588 bastu 1
7589 basunstöt 3
7590 basvattenförbrukning 1
7591 baxa 1
7592 bayerska 1
7593 bayerskt 1
7594 bayrare 1
7595 be 63
7596 beakta 29
7597 beaktades 5
7598 beaktande 7
7599 beaktanden 1
7600 beaktandet 2
7601 beaktansvärt 1
7602 beaktar 13
7603 beaktas 29
7604 beaktat 8
7605 beaktats 7
7606 bearbeta 2
7607 bearbetade 1
7608 bearbetande 1
7609 bearbetas 1
7610 beblandade 1
7611 bebodd 1
7612 bebodda 2
7613 bebyggelse 1
7614 bebyggelsen 1
7615 bebådade 1
7616 bedra 3
7617 bedragare 1
7618 bedrar 2
7619 bedrevs 1
7620 bedrifter 1
7621 bedriva 15
7622 bedrivas 5
7623 bedriver 12
7624 bedrivit 3
7625 bedrivs 6
7626 bedrägeri 15
7627 bedrägeribekämpning 7
7628 bedrägeribekämpningen 1
7629 bedrägerier 15
7630 bedrägerierna 1
7631 bedrägeriet 2
7632 bedrägerikonventionen 1
7633 bedrägerimål 1
7634 bedräglig 1
7635 bedrövelser 1
7636 bedrövliga 1
7637 bedrövligt 2
7638 bedöma 29
7639 bedömas 8
7640 bedömda 1
7641 bedömdes 1
7642 bedömer 11
7643 bedömning 41
7644 bedömningar 4
7645 bedömningarna 2
7646 bedömningen 8
7647 bedöms 8
7648 bedömt 2
7649 beef 1
7650 befallningar 1
7651 befann 9
7652 befara 2
7653 befarar 5
7654 befatta 2
7655 befattar 1
7656 befattat 4
7657 befattning 3
7658 befattningar 4
7659 befattningarna 1
7660 befinna 9
7661 befinner 92
7662 befintlig 2
7663 befintliga 49
7664 befintligt 1
7665 befläckad 1
7666 befogad 3
7667 befogade 3
7668 befogat 4
7669 befogenhet 11
7670 befogenheter 45
7671 befogenheterna 2
7672 befogenhetsområden 1
7673 befolka 1
7674 befolkad 1
7675 befolkade 6
7676 befolkning 34
7677 befolkningar 4
7678 befolkningarna 10
7679 befolkningarnas 2
7680 befolkningen 87
7681 befolkningens 10
7682 befolknings 1
7683 befolkningsdelar 1
7684 befolkningsgrupper 10
7685 befolkningsgrupperna 4
7686 befolkningskoncentration 1
7687 befolkningslager 1
7688 befolkningslagren 1
7689 befolkningsmajoriteten 2
7690 befolkningsmajoritetens 1
7691 befolkningssammansättningen 1
7692 befolkningssiffra 2
7693 befolkningsspridning 1
7694 befolkningsstorlek 1
7695 befolkningsstorleken 1
7696 befolkningsstruktur 1
7697 befolkningstillväxt 1
7698 befolkningstäthet 1
7699 befolkningstätheten 1
7700 befolkningsunderlag 1
7701 befordran 7
7702 befordras 1
7703 befraktare 1
7704 befraktaren 4
7705 befraktarna 2
7706 befraktarnas 3
7707 befria 1
7708 befriad 2
7709 befriar 1
7710 befrias 5
7711 befriat 1
7712 befriats 1
7713 befrukta 1
7714 befrämjandet 1
7715 befrämjat 1
7716 befullmäktigade 1
7717 befunnit 3
7718 befunnits 1
7719 befäl 2
7720 befälet 2
7721 befälhavare 2
7722 befälhavaren 1
7723 befängda 2
7724 befängt 1
7725 befäst 1
7726 befästa 11
7727 befästande 1
7728 befäste 1
7729 befäster 3
7730 befästes 1
7731 begagnade 6
7732 begav 1
7733 bege 3
7734 begrava 1
7735 begravning 3
7736 begravningsplatser 1
7737 begrep 2
7738 begrepp 17
7739 begreppen 5
7740 begreppet 31
7741 begripa 2
7742 begriper 4
7743 begriplig 1
7744 begripligare 1
7745 begripligt 3
7746 begrunda 3
7747 begrundade 1
7748 begränsa 41
7749 begränsad 37
7750 begränsade 27
7751 begränsades 2
7752 begränsande 2
7753 begränsar 19
7754 begränsas 17
7755 begränsat 15
7756 begränsats 1
7757 begränsning 11
7758 begränsningar 20
7759 begränsningarna 6
7760 begränsningen 1
7761 begränsningsavtal 1
7762 begynnande 1
7763 begynnelsebokstaven 1
7764 begynnelsen 2
7765 begynte 1
7766 begär 42
7767 begära 21
7768 begäran 63
7769 begäran.)Beträffande 1
7770 begäras 3
7771 begärda 1
7772 begärde 12
7773 begärets 1
7774 begärs 8
7775 begärt 24
7776 begå 3
7777 begångna 1
7778 begår 3
7779 begås 6
7780 begått 5
7781 begåtts 3
7782 begåvning 1
7783 behag 1
7784 behagligt 1
7785 behandla 36
7786 behandlad 1
7787 behandlade 5
7788 behandlades 6
7789 behandlar 38
7790 behandlas 49
7791 behandlat 10
7792 behandlats 4
7793 behandling 35
7794 behandlingarna 1
7795 behandlingen 48
7796 behandlingens 1
7797 behandlingsanläggning 1
7798 behandlingsanläggningarna 1
7799 behandlingscentraler 1
7800 behov 86
7801 behoven 12
7802 behovet 97
7803 behäftat 1
7804 behärskade 1
7805 behåll 1
7806 behålla 33
7807 behållare 1
7808 behållas 1
7809 behåller 2
7810 behållit 1
7811 behållits 1
7812 behålls 1
7813 behöll 3
7814 behölls 1
7815 behörig 2
7816 behöriga 15
7817 behörige 1
7818 behörighet 16
7819 behörigheten 2
7820 behörigheter 4
7821 behörighetsnivå 1
7822 behörighetsområde 4
7823 behörighetsområden 1
7824 behörigt 1
7825 behöva 50
7826 behövande 1
7827 behövas 6
7828 behövde 10
7829 behövdes 3
7830 behöver 264
7831 behövliga 1
7832 behövs 113
7833 behövt 3
7834 behövts 1
7835 beivras 1
7836 bekant 10
7837 bekanta 3
7838 bekantgjorts 1
7839 beklaga 20
7840 beklagade 2
7841 beklagande 6
7842 beklaganden 3
7843 beklagansvärd 1
7844 beklagansvärda 2
7845 beklagansvärt 3
7846 beklagar 49
7847 beklagat 2
7848 beklaglig 2
7849 beklagliga 3
7850 beklagligt 17
7851 beklämmande 2
7852 bekom 1
7853 bekostat 1
7854 bekostnad 7
7855 bekräfta 39
7856 bekräftade 5
7857 bekräftades 3
7858 bekräftande 1
7859 bekräftar 17
7860 bekräftas 9
7861 bekräftat 7
7862 bekräftats 4
7863 bekräftelse 5
7864 bekräftelsen 2
7865 bekväm 1
7866 bekvämligheter 2
7867 bekvämlighetsflagg 23
7868 bekvämlighetsflaggade 5
7869 bekvämlighetsflaggades 1
7870 bekvämlighetsflaggen 1
7871 bekvämlighetsflaggningen 1
7872 bekvämt 3
7873 bekymmer 17
7874 bekymmersamma 1
7875 bekymmersamt 3
7876 bekymra 1
7877 bekymrad 9
7878 bekymrade 8
7879 bekymrande 1
7880 bekymrar 7
7881 bekymrat 2
7882 bekämpa 76
7883 bekämpade 2
7884 bekämpande 3
7885 bekämpandet 2
7886 bekämpar 6
7887 bekämpas 3
7888 bekämpats 1
7889 bekämpning 13
7890 bekämpningen 5
7891 bekämpningsmedel 1
7892 bekänna 1
7893 bekännelse 1
7894 bekännelser 1
7895 bekänner 1
7896 belagda 1
7897 belagt 1
7898 belasta 1
7899 belastande 1
7900 belastar 2
7901 belastas 2
7902 belastning 4
7903 belastningar 1
7904 belgisk 3
7905 belgiska 13
7906 belopp 15
7907 beloppen 3
7908 beloppet 6
7909 beloppets 1
7910 belysa 2
7911 belysas 1
7912 belyser 2
7913 belysning 2
7914 belyst 2
7915 beläget 2
7916 belägg 1
7917 beläggs 1
7918 belägna 7
7919 belåtenhet 2
7920 belåtet 3
7921 belåtna 1
7922 belönar 1
7923 belönas 2
7924 belöpte 1
7925 bemanningsbehovet 1
7926 bemyndigande 6
7927 bemyndigar 1
7928 bemärkelse 4
7929 bemärkelsen 4
7930 bemästra 1
7931 bemöda 5
7932 bemödanden 4
7933 bemödar 1
7934 bemöta 10
7935 bemötande 1
7936 bemötas 1
7937 bemöter 5
7938 bemöts 2
7939 bemötts 1
7940 ben 10
7941 bench-marking 1
7942 benchmark 1
7943 benchmarking 3
7944 benchmarking-system 1
7945 benchmarks 1
7946 benen 4
7947 benet 1
7948 benhård 1
7949 benhårda 1
7950 benhårt 1
7951 benig 1
7952 benmjöl 1
7953 bensin 2
7954 bensinpriset 1
7955 benstomme 2
7956 benägna 3
7957 benämning 1
7958 benämns 1
7959 benåda 1
7960 beordra 1
7961 beordrat 1
7962 beordrats 1
7963 ber 101
7964 bereda 2
7965 beredas 1
7966 beredd 46
7967 beredda 44
7968 bereder 1
7969 beredningen 1
7970 bereds 1
7971 beredskap 3
7972 beredskapen 1
7973 beredvilligt 1
7974 berett 8
7975 beretts 2
7976 berg 5
7977 berget 2
7978 bergs- 1
7979 bergskommunerna 1
7980 bergsområden 1
7981 bergssektorer 1
7982 bergssidan 1
7983 berika 7
7984 berikande 2
7985 berikar 3
7986 berikas 1
7987 berikat 1
7988 bero 1
7989 berodde 6
7990 beroende 63
7991 beroendeminskning 1
7992 beroendet 3
7993 beror 54
7994 berott 2
7995 berusa 1
7996 berusad 2
7997 berusat 1
7998 beryktad 1
7999 beryktade 1
8000 beräkna 4
8001 beräknade 3
8002 beräknades 1
8003 beräknar 2
8004 beräknas 6
8005 beräknat 2
8006 beräknats 1
8007 beräkning 2
8008 beräkningar 4
8009 beräkningarna 4
8010 beräkningen 8
8011 berätta 24
8012 berättade 16
8013 berättar 5
8014 berättare 1
8015 berättas 1
8016 berättat 4
8017 berättelse 4
8018 berättelsen 2
8019 berättelserna 1
8020 berättiga 1
8021 berättigad 9
8022 berättigade 18
8023 berättigande 6
8024 berättigar 3
8025 berättigas 2
8026 berättigat 13
8027 berömd 2
8028 berömda 6
8029 berömde 1
8030 berömma 5
8031 berömmande 1
8032 berömt 1
8033 berömvärd 1
8034 berömvärda 2
8035 berömvärt 2
8036 berör 43
8037 beröra 2
8038 beröras 4
8039 berörd 2
8040 berörda 62
8041 berörde 4
8042 berördes 2
8043 beröring 1
8044 beröringen 1
8045 beröringspunkter 1
8046 berörs 21
8047 berört 8
8048 berörts 3
8049 beröva 3
8050 berövar 1
8051 berövats 1
8052 besatta 1
8053 besatthet 1
8054 besegla 1
8055 besegrade 1
8056 besegrades 1
8057 besegrar 1
8058 besiktning 1
8059 besiktningar 1
8060 besiktningsinstrument 1
8061 besiktningsmyndigheterna 1
8062 besitter 5
8063 beskaffenhet 1
8064 beskatta 2
8065 beskattad 1
8066 beskattas 1
8067 beskattning 9
8068 beskattningen 2
8069 beskattningsfrågor 1
8070 beskattningskod 1
8071 besked 12
8072 beskjuta 1
8073 beskrev 5
8074 beskrevs 2
8075 beskriva 9
8076 beskrivande 2
8077 beskrivas 3
8078 beskriver 7
8079 beskrivet 2
8080 beskrivit 9
8081 beskrivits 2
8082 beskrivna 2
8083 beskrivning 12
8084 beskrivningar 1
8085 beskrivs 10
8086 beskydd 6
8087 beskydda 1
8088 beskylla 1
8089 beskyller 1
8090 beskyllningar 1
8091 beskylls 1
8092 beskyllts 1
8093 beskåda 1
8094 besköt 1
8095 beslag 1
8096 beslagta 1
8097 beslagtagna 1
8098 beslut 264
8099 besluta 27
8100 beslutade 22
8101 beslutades 5
8102 beslutande 2
8103 beslutandefrihet 1
8104 beslutandemakten 1
8105 beslutandeplanet 1
8106 beslutanderätt 2
8107 beslutar 13
8108 beslutas 8
8109 beslutat 15
8110 beslutats 6
8111 besluten 29
8112 beslutet 38
8113 beslutets 1
8114 beslutna 3
8115 besluts- 2
8116 beslutsam 4
8117 beslutsamhet 17
8118 beslutsamma 1
8119 beslutsamt 10
8120 beslutscentrum 2
8121 beslutscentrumen 1
8122 beslutsfattande 22
8123 beslutsfattandet 10
8124 beslutsfattandets 1
8125 beslutsfattare 5
8126 beslutsfattarna 5
8127 beslutsfrihet 1
8128 beslutsförfaranden 1
8129 beslutsförfarandena 1
8130 beslutsförfarandet 1
8131 beslutsmakt 1
8132 beslutsmakten 2
8133 beslutsnivå 1
8134 beslutsorgan 1
8135 beslutsposter 1
8136 beslutsprocess 4
8137 beslutsprocessen 25
8138 beslutsprocesser 2
8139 beslutsprocesserna 4
8140 beslutsrätt 3
8141 beslutsstrukturer 1
8142 beslutstyperna 1
8143 beslutsunderlag 1
8144 beslutsunderlaget 2
8145 besläktade 1
8146 beslöt 13
8147 bespara 3
8148 besparade 1
8149 besparar 2
8150 besparingar 6
8151 besparings- 1
8152 best 4
8153 bestod 6
8154 bestraffa 1
8155 bestraffade 1
8156 bestraffar 2
8157 bestraffas 6
8158 bestraffning 1
8159 bestraffningar 1
8160 bestrida 4
8161 bestrider 1
8162 bestrids 2
8163 bestrålning 1
8164 bestyrka 1
8165 beställa 1
8166 beställde 2
8167 beställdes 1
8168 beställningar 1
8169 beställt 2
8170 beställts 1
8171 bestämd 7
8172 bestämda 13
8173 bestämdaste 2
8174 bestämde 4
8175 bestämdhet 2
8176 bestämma 22
8177 bestämmas 2
8178 bestämmelse 11
8179 bestämmelsen 3
8180 bestämmelsens 1
8181 bestämmelser 114
8182 bestämmelserna 56
8183 bestämmer 8
8184 bestäms 4
8185 bestämt 40
8186 bestämts 1
8187 beständig 2
8188 bestå 8
8189 bestående 14
8190 bestånd 8
8191 bestånden 8
8192 beståndet 3
8193 beståndsdel 11
8194 beståndsdelar 15
8195 beståndsdelarna 3
8196 beståndsdelen 1
8197 består 41
8198 bestått 1
8199 bestört 1
8200 bestörtning 3
8201 besvara 30
8202 besvarade 2
8203 besvarades 1
8204 besvarandet 1
8205 besvarar 4
8206 besvaras 9
8207 besvarat 1
8208 besvarats 2
8209 besvikelse 9
8210 besviken 8
8211 besviket 1
8212 besvikna 5
8213 besvär 2
8214 besvära 1
8215 besvärades 1
8216 besväret 3
8217 besvärlig 5
8218 besvärliga 5
8219 besvärligare 2
8220 besvärligt 2
8221 besynnerlig 2
8222 besynnerliga 2
8223 besynnerligheter 2
8224 besynnerligt 1
8225 besättning 3
8226 besättningen 2
8227 besök 27
8228 besöka 7
8229 besökare 1
8230 besöket 2
8231 besöksnäringens 1
8232 besökte 5
8233 beta 1
8234 betade 1
8235 betala 83
8236 betalade 4
8237 betalar 48
8238 betalas 6
8239 betalat 6
8240 betalats 7
8241 betalbara 1
8242 betalbart 1
8243 betald 1
8244 betalda 2
8245 betalning 2
8246 betalningar 6
8247 betalningen 1
8248 betalningsansvariga 1
8249 betalningsbemyndiganden 1
8250 betalningsförmågan 1
8251 betalningsförseningar 1
8252 betalningsmedel 1
8253 betalningsskyldiges 1
8254 betalningssystemen 1
8255 betalt 5
8256 betalts 1
8257 bete 1
8258 beteckna 3
8259 betecknade 1
8260 betecknande 2
8261 betecknar 2
8262 betecknas 5
8263 beteckningen 3
8264 beteende 4
8265 beteendemönster 1
8266 beteenden 1
8267 beter 1
8268 betingad 1
8269 betingade 1
8270 betingar 1
8271 betingat 1
8272 betingelser 3
8273 betingelserna 1
8274 betitlat 1
8275 betjäna 3
8276 betjänas 1
8277 betjänta 1
8278 betona 67
8279 betonade 11
8280 betonades 2
8281 betonandet 1
8282 betonar 27
8283 betonas 18
8284 betonat 10
8285 betonats 1
8286 betoning 5
8287 betoningen 1
8288 betrakta 18
8289 betraktade 6
8290 betraktande 2
8291 betraktar 26
8292 betraktas 25
8293 betraktat 3
8294 betraktats 1
8295 betryggande 5
8296 beträda 1
8297 beträffade 1
8298 beträffande 68
8299 beträffar 94
8300 bett 12
8301 betungande 3
8302 betvivla 2
8303 betvivlade 1
8304 betvivlar 9
8305 betyda 7
8306 betydande 68
8307 betydde 6
8308 betydelse 146
8309 betydelsefull 11
8310 betydelsefulla 16
8311 betydelsefullt 17
8312 betydelselös 1
8313 betydelselöst 2
8314 betydelsen 28
8315 betyder 60
8316 betydligt 32
8317 betyg 1
8318 betygar 1
8319 betänk 1
8320 betänka 5
8321 betänkande 380
8322 betänkanden 25
8323 betänkandena 5
8324 betänkandet 198
8325 betänkandets 4
8326 betänker 3
8327 betänkligheter 7
8328 beundran 1
8329 beundrar 4
8330 beundrat 1
8331 bevaka 5
8332 bevakad 1
8333 bevakade 1
8334 bevakar 3
8335 bevakaren 1
8336 bevakning 2
8337 bevara 54
8338 bevarad 2
8339 bevarande 26
8340 bevarandeområde 2
8341 bevarandet 12
8342 bevarar 5
8343 bevaras 6
8344 bevarats 2
8345 bevattning 3
8346 beveka 1
8347 bevekande 1
8348 bevilja 24
8349 beviljad 1
8350 beviljade 6
8351 beviljades 1
8352 beviljande 4
8353 beviljanden 2
8354 beviljandet 4
8355 beviljar 9
8356 beviljas 12
8357 beviljat 7
8358 beviljats 8
8359 bevis 50
8360 bevisa 11
8361 bevisad 1
8362 bevisade 1
8363 bevisades 1
8364 bevisar 3
8365 bevisas 1
8366 bevisat 2
8367 bevisats 3
8368 bevisbörda 3
8369 bevisbördan 5
8370 bevisen 4
8371 beviset 3
8372 bevisningsfel 1
8373 bevista 1
8374 bevistade 1
8375 bevittna 2
8376 bevittnar 3
8377 bevittnat 2
8378 bevänt 1
8379 beväpning 1
8380 bibehålla 19
8381 bibehållande 1
8382 bibehållandet 1
8383 bibehållas 3
8384 bibehållen 2
8385 bibehåller 5
8386 bibehållits 1
8387 bibehålls 4
8388 biblioteken 1
8389 bibliotekens 1
8390 bidade 1
8391 bidra 103
8392 bidrag 102
8393 bidragande 2
8394 bidragen 7
8395 bidraget 7
8396 bidragit 19
8397 bidragsberoende 1
8398 bidragsgivare 3
8399 bidragsgivaren 3
8400 bidragsgivarna 4
8401 bidragsgivning 1
8402 bidragshjälp 1
8403 bidragsnarkomaner 1
8404 bidrar 52
8405 bidrog 6
8406 bieffekt 1
8407 bieffekter 2
8408 bieffekterna 1
8409 bifall 7
8410 bifalla 1
8411 bifallas 3
8412 bifallit 1
8413 biff 1
8414 bifloder 1
8415 bifogade 1
8416 bifogat 1
8417 bifångster 1
8418 bifångsterna 1
8419 biföll 4
8420 big 1
8421 bigotteri 1
8422 bil 19
8423 bil- 1
8424 bilaga 6
8425 bilagan 3
8426 bilagor 1
8427 bilagorna 3
8428 bilagts 1
8429 bilar 62
8430 bilarbetare 1
8431 bilarna 8
8432 bilarnas 2
8433 bilatera 1
8434 bilateral 3
8435 bilaterala 12
8436 bilateralt 6
8437 bilbeståndet 1
8438 bilbranschen 1
8439 bild 34
8440 bilda 14
8441 bildade 2
8442 bildades 4
8443 bildande 2
8444 bildandet 8
8445 bildar 10
8446 bildas 11
8447 bildat 2
8448 bildats 2
8449 bildelar 2
8450 bildelarna 1
8451 bilden 9
8452 bilder 3
8453 bilderna 1
8454 bildligt 1
8455 bildningar 1
8456 bildnings- 1
8457 bildtext 1
8458 bilen 22
8459 bilens 1
8460 bilindustri 6
8461 bilindustrin 18
8462 bilindustrins 5
8463 bilindustris 2
8464 bilister 1
8465 bilisterna 1
8466 biljetten 1
8467 biljoner 1
8468 bilkonstruktörerna 1
8469 bilkyrkogårdar 1
8470 bilköpare 2
8471 billig 1
8472 billiga 2
8473 billigare 6
8474 billigaste 1
8475 billigt 4
8476 bilmärke 1
8477 bilolyckan 1
8478 bilpark 2
8479 bilparken 4
8480 bilpriset 1
8481 bilproduktion 1
8482 bils 2
8483 bilsektorns 1
8484 bilskrotningen 1
8485 bilskrotningsmetod 1
8486 biltillverkare 4
8487 biltillverkaren 1
8488 biltillverkares 1
8489 biltillverkarna 8
8490 biltillverkarnas 1
8491 biltillverkning 1
8492 bilvrak 4
8493 bilvraket 2
8494 bilägarna 1
8495 bilägga 1
8496 bilåtervinningsmarknaden 1
8497 bin 2
8498 binda 4
8499 bindande 34
8500 bindas 1
8501 binder 3
8502 bio 2
8503 biodiversitet 1
8504 biografi 1
8505 biologer 1
8506 biologisk 8
8507 biologiska 22
8508 biologiskt 2
8509 biomassa 1
8510 bioplast 1
8511 biosfären 1
8512 biosäkerhet 1
8513 biosäkerhetsprotokollet 1
8514 biotekniken 2
8515 biotekniska 1
8516 biotoperna 1
8517 bisarra 1
8518 bister 1
8519 bistå 7
8520 bistånd 41
8521 biståndet 10
8522 bistånds 1
8523 biståndsflödena 2
8524 biståndsfrågor 1
8525 biståndsgivare 1
8526 biståndsgivaren 4
8527 biståndshjälp 1
8528 biståndsideologin 1
8529 biståndsmottagare 1
8530 biståndspengarna 2
8531 biståndspolitik 1
8532 biståndspolitiken 1
8533 biståndsprogram 1
8534 biståndsprogrammen 2
8535 biståndssystem 1
8536 biståndsvolym 1
8537 bistår 1
8538 bistått 3
8539 bit 10
8540 bitande 1
8541 bitar 3
8542 biter 2
8543 bitmappar 1
8544 biträdande 1
8545 biträdas 1
8546 biträde 1
8547 bitter 3
8548 bitterhet 1
8549 bittert 1
8550 bittra 1
8551 bjuda 5
8552 bjudande 1
8553 bjuder 2
8554 bjudit 2
8555 bjärt 1
8556 bjärtare 1
8557 bjöd 2
8558 bl 3
8559 bl.a. 49
8560 blackmail 1
8561 blad 1
8562 bladen 1
8563 blamerande 1
8564 bland 158
8565 blanda 11
8566 blandad 1
8567 blandade 2
8568 blandar 4
8569 blandas 4
8570 blandat 2
8571 blandning 5
8572 blandningar 1
8573 blandningen 1
8574 blandningens 1
8575 blandskogar 1
8576 blanka 1
8577 blanketter 1
8578 blanko 1
8579 blanksteg 1
8580 blankt 1
8581 bleckhink 1
8582 bleiben 1
8583 blek 1
8584 bleka 5
8585 blekaste 1
8586 blekgult 1
8587 bleknat 1
8588 blekningsmedel 1
8589 blekt 1
8590 blev 99
8591 bli 413
8592 blick 10
8593 blicka 1
8594 blickar 4
8595 blickarna 1
8596 blicken 8
8597 blickfältet 1
8598 blickpunkten 1
8599 blind 4
8600 blinda 2
8601 blinkade 3
8602 blint 4
8603 blir 305
8604 blivande 1
8605 blivit 103
8606 blixt 2
8607 blixtar 1
8608 blixtlås 1
8609 blixtrande 1
8610 blixtvisit 1
8611 blixtärr 1
8612 block 3
8613 blockad 3
8614 blockaden 7
8615 blockadinstrument 1
8616 blockbildning 1
8617 blockera 5
8618 blockerad 2
8619 blockerade 2
8620 blockerar 4
8621 blockeras 3
8622 blockerat 3
8623 blockering 1
8624 blocket 1
8625 blod 6
8626 blodbad 1
8627 blodet 1
8628 blodfläckad 1
8629 blodigt 2
8630 blodspillan 1
8631 blomma 2
8632 blommig 1
8633 blommiga 1
8634 blommigt 1
8635 blommor 4
8636 blomrabatterna 1
8637 blomsternoter 1
8638 blomstrande 1
8639 blomstrar 1
8640 blomstring 2
8641 blond 3
8642 blonda 1
8643 blonde 1
8644 blott 2
8645 blotta 1
8646 blottade 1
8647 blottades 1
8648 blottas 1
8649 blunda 4
8650 blundar 4
8651 bly 5
8652 blyga 1
8653 blyghet 1
8654 blygrått 1
8655 blygsam 3
8656 blygsamhet 2
8657 blygsamma 6
8658 blygsammare 1
8659 blygsamt 1
8660 blyregnet 1
8661 bländande 4
8662 blänka 1
8663 blänkande 1
8664 blänkte 2
8665 blå 11
8666 blåa 1
8667 blåfenad 8
8668 blåfenade 3
8669 blågrön 1
8670 blåkläder 1
8671 blåsa 1
8672 blåser 1
8673 blåslagen 1
8674 blåste 3
8675 blått 2
8676 blöt 2
8677 bo 8
8678 bodde 10
8679 boende 3
8680 bogsera 2
8681 bogserade 1
8682 bogserarna 1
8683 bogserbåt 2
8684 bogserbåtar 1
8685 bojkott 1
8686 bojkotta 1
8687 bojkottar 1
8688 bojkotten 1
8689 bok 15
8690 bokad 1
8691 boken 4
8692 bokens 1
8693 bokföringsbegrepp 1
8694 bokhandeln 2
8695 boklista 1
8696 bokmärket 1
8697 bokslut 3
8698 bokstaven 1
8699 bokstavligen 5
8700 bokstavligt 1
8701 bokälskare 1
8702 bolag 7
8703 bolagen 2
8704 bolagens 2
8705 bolaget 4
8706 bolagets 1
8707 bolags 2
8708 bolagsskatter 2
8709 bollen 3
8710 bolsjevikiska 1
8711 bolsjevitisk 1
8712 bomb 7
8713 bomba 1
8714 bombades 1
8715 bombarderade 1
8716 bombattentat 1
8717 bomben 1
8718 bomber 2
8719 bombexplosioner 1
8720 bombning 1
8721 bombningar 6
8722 bombningarna 5
8723 bombningen 1
8724 bomull 1
8725 bomullstyger 1
8726 bon 1
8727 bondens 1
8728 bondgård 1
8729 bondgården 1
8730 bondkvinna 1
8731 bonus 1
8732 booming 1
8733 bor 44
8734 bord 10
8735 borde 237
8736 bordeauxvin 1
8737 borden 1
8738 bordet 9
8739 bordlades 1
8740 bords 1
8741 bordsgaffeln 1
8742 bordsgrannens 1
8743 borga 1
8744 borgar 2
8745 borgen 1
8746 borgenärernas 1
8747 borgerlig 1
8748 borgmästare 8
8749 borgmästarens 1
8750 borgmästarinna 1
8751 borgmästarna 1
8752 borrar 3
8753 borsta 2
8754 borstade 1
8755 bort 127
8756 borta 10
8757 bortemot 1
8758 bortfaller 8
8759 bortfallet 2
8760 bortförd 1
8761 bortglömd 2
8762 bortglömda 2
8763 bortkastad 1
8764 bortkastat 2
8765 bortom 15
8766 bortprioriteras 1
8767 bortse 11
8768 bortser 6
8769 bortsett 8
8770 bortskämda 2
8771 bortsållningen 1
8772 borttagandet 1
8773 borttappat 1
8774 bortåt 1
8775 bosatt 1
8776 bosatta 6
8777 boskapsdöden 1
8778 boskapsinitiativ 1
8779 boskapsskötarnas 1
8780 boskapsskötsel 2
8781 boskapsuppfödarna 1
8782 bosnier 2
8783 bostad 1
8784 bostaden 1
8785 bostadshyror 1
8786 bostadsprojekt 1
8787 bostäder 7
8788 bosätta 3
8789 bosättare 1
8790 bosättningar 5
8791 bosättningarna 7
8792 bosättningsdirektiven 1
8793 bosättningsområdena 1
8794 bosättningsvillkoren 1
8795 bot 3
8796 bota 1
8797 botade 1
8798 botar 2
8799 botemedlet 2
8800 bott 2
8801 botten 19
8802 bottenlös 1
8803 bottenlösa 1
8804 bottnar 3
8805 bottnen 1
8806 bottom-up-koncept 1
8807 bovar 1
8808 boven 2
8809 boy 1
8810 bra 272
8811 bragdes 1
8812 brakade 1
8813 brand 2
8814 branden 1
8815 brandgula 1
8816 brandmän 1
8817 brann 1
8818 bransch 5
8819 branschen 5
8820 branscher 3
8821 branscherna 3
8822 brant 1
8823 branten 2
8824 brasan 3
8825 brast 4
8826 brave 1
8827 bred 21
8828 breda 17
8829 bredare 22
8830 bredast 2
8831 bredband 1
8832 bredbandsnät 1
8833 bredda 5
8834 breddar 1
8835 bredde 2
8836 bredden 4
8837 breddgraden 1
8838 breder 1
8839 bredvid 14
8840 bretagniska 1
8841 bretonne 1
8842 bretonska 3
8843 brett 20
8844 brev 29
8845 brevbärare 1
8846 brevbäraren 7
8847 brevbärarens 1
8848 brevet 3
8849 brevinsamling 1
8850 brevlåda 1
8851 brevlådeföretag 1
8852 brevutbärning 1
8853 brevväxlingen 1
8854 bricka 1
8855 brickan 2
8856 brickorna 2
8857 briefing-PM 1
8858 brigad 1
8859 briljera 1
8860 brillorna 1
8861 bringa 6
8862 bringan 1
8863 bringar 1
8864 bringas 1
8865 bringat 1
8866 brinna 1
8867 brinnande 1
8868 brinner 1
8869 bris 1
8870 briserande 1
8871 briserat 1
8872 brist 55
8873 brista 1
8874 bristande 24
8875 bristen 42
8876 brister 42
8877 bristerna 10
8878 bristfällig 5
8879 bristfälliga 6
8880 bristfälligt 4
8881 brits 1
8882 britter 2
8883 brittisk 4
8884 brittiska 36
8885 brittiske 1
8886 brittiskt 4
8887 bro 4
8888 broar 4
8889 broderade 1
8890 broders 1
8891 broderskap 4
8892 broförbindelse 1
8893 brohuvuden 1
8894 brokig 1
8895 brokigt 1
8896 bromerade 5
8897 broms 1
8898 bromsa 5
8899 bromsar 4
8900 bromsas 1
8901 bromsat 1
8902 bromsen 1
8903 bromsvätska 1
8904 bronsmynten 1
8905 bror 2
8906 broregioner 1
8907 brorsdotter 1
8908 broskbemängda 1
8909 brother 1
8910 brott 54
8911 brottas 2
8912 brottats 2
8913 brotten 2
8914 brottmål 15
8915 brottmålsdomstol 1
8916 brottmålsdomstolar 1
8917 brottmålsdomstolen 3
8918 brottningsmatchen 1
8919 brottsanklagar 1
8920 brottsbekämpning 3
8921 brottsbekämpningen 2
8922 brottsfrågor 1
8923 brottsförebyggande 1
8924 brottslig 1
8925 brottsliga 4
8926 brottslighet 9
8927 brottsligheten 15
8928 brottsling 1
8929 brottslingar 3
8930 brottslingarna 2
8931 brottsmålssidan 1
8932 brottsoffer 2
8933 brottsrubriker 1
8934 brottsskolor 1
8935 brotullarna 1
8936 bruk 14
8937 brukade 24
8938 brukar 8
8939 brukarna 1
8940 brukas 1
8941 bruket 7
8942 brummade 2
8943 brun 1
8944 bruna 4
8945 brunn 1
8946 brunnen 1
8947 brunrosa 1
8948 brusande 1
8949 bruset 1
8950 brutal 1
8951 brutala 4
8952 brutalt 2
8953 brutit 5
8954 brutits 3
8955 bruttoinvesteringar 1
8956 bruttonationalinkomsten 3
8957 bruttonationalprodukt 2
8958 bruttonationalprodukten 2
8959 bry 5
8960 brydde 4
8961 brygga 1
8962 bryggan 1
8963 brynet 1
8964 bryr 12
8965 brysk 1
8966 bryta 16
8967 brytas 2
8968 bryter 18
8969 brytning 4
8970 brytningar 1
8971 brytningen 2
8972 brytningsåret 1
8973 bryts 1
8974 brytt 1
8975 bräcklig 2
8976 bräckliga 4
8977 bräm 1
8978 brända 2
8979 brände 2
8980 bränder 1
8981 bränderna 1
8982 bränna 3
8983 brännande 1
8984 brännas 1
8985 bränning 2
8986 bränningar 1
8987 bränningarna 1
8988 bränningen 1
8989 brännmärka 1
8990 bränsle 3
8991 bränsleförvaring 1
8992 bränslekvaliteten 1
8993 bränslen 3
8994 bränsleskatt 1
8995 bränslesnåla 2
8996 bränslesnålare 2
8997 bränslet 1
8998 bränsletransporter 1
8999 bränts 1
9000 bräsch 1
9001 bräschen 2
9002 brådska 4
9003 brådskande 44
9004 brådskar 2
9005 bråk 1
9006 bråkdel 2
9007 bråkdels 1
9008 bråket 1
9009 bråkiga 1
9010 bröd 6
9011 bröder 1
9012 brödskiva 1
9013 brödsäd 1
9014 bröllopsnatten 1
9015 bröst 4
9016 brösten 2
9017 bröstet 1
9018 brösttoner 1
9019 bröt 6
9020 bubbla 1
9021 bubblan 2
9022 bubblor 1
9023 bucklade 1
9024 buddha 1
9025 buddhistiska 1
9026 budfirmor 1
9027 budget 52
9028 budgetanslag 4
9029 budgetanslaget 1
9030 budgetanspråk 1
9031 budgetar 6
9032 budgetarbetet 1
9033 budgetarna 1
9034 budgetbalans 1
9035 budgetbehov 1
9036 budgetbeloppet 1
9037 budgetberäkning 1
9038 budgetberäkningen 1
9039 budgetbeslut 1
9040 budgetbestämmelserna 1
9041 budgetchefen 1
9042 budgetdiskussioner 1
9043 budgeteffekten 1
9044 budgeten 53
9045 budgetenhet 1
9046 budgetens 1
9047 budgetera 1
9048 budgetfråga 1
9049 budgetfrågan 3
9050 budgetfrågor 1
9051 budgetförfarande 1
9052 budgetförfarandet 2
9053 budgetförordning 2
9054 budgetförordningen 8
9055 budgetförslag 1
9056 budgetförslaget 2
9057 budgetförvaltning 2
9058 budgetgest 1
9059 budgetkonsekvenser 2
9060 budgetkontroll 1
9061 budgetkontrollen 1
9062 budgetkontrollutskott 1
9063 budgetkontrollutskottet 14
9064 budgetkontrollutskottets 1
9065 budgetkravet 1
9066 budgetmyndigheten 2
9067 budgetmässiga 2
9068 budgetnivå 1
9069 budgetnärmanden 1
9070 budgetområde 1
9071 budgetplan 6
9072 budgetplanen 9
9073 budgetplaner 1
9074 budgetplanerna 3
9075 budgetpolitik 5
9076 budgetpolitiken 1
9077 budgetpost 13
9078 budgetposten 7
9079 budgetposter 5
9080 budgetposterna 2
9081 budgetreform 1
9082 budgetrubrik 3
9083 budgetrubriker 1
9084 budgetsituation 1
9085 budgetstöd 1
9086 budgetstödet 1
9087 budgetsynpunkt 1
9088 budgetunderskott 1
9089 budgetutskott 1
9090 budgetutskottet 10
9091 budgetåret 13
9092 budgetårets 1
9093 budgetåtgärder 1
9094 budgetöverbud 1
9095 budgetöverenskommelse 1
9096 budgetövervakare 1
9097 budord 1
9098 budordet 1
9099 buds 2
9100 budskap 23
9101 budskapet 5
9102 bugade 1
9103 building 1
9104 buk 1
9105 bukiga 1
9106 bukt 2
9107 bukter 1
9108 bullar 2
9109 bulldozrar 1
9110 bulle 1
9111 buller 1
9112 bullrigare 1
9113 bultade 1
9114 bunden 3
9115 bundna 1
9116 bundsförvant 1
9117 bur 5
9118 burden 1
9119 buren 2
9120 burens 1
9121 burit 6
9122 burken 1
9123 burklocket 1
9124 burktomater 1
9125 busflin 1
9126 bushen 3
9127 business 1
9128 business-toppmötet 1
9129 buskagen 1
9130 buskiga 1
9131 buskvegetationen 1
9132 buss 4
9133 bussar 2
9134 bussfilerna 1
9135 busslinjer 1
9136 busstjänst 1
9137 but 1
9138 butelj 1
9139 butik 2
9140 butiken 4
9141 butiker 2
9142 butiksdörren 1
9143 butiksfönster 1
9144 butiksfönstren 1
9145 butiksfönstret 1
9146 butiksförsäljningen 1
9147 buttert 1
9148 buxbomsbord 1
9149 bwana 1
9150 by 6
9151 byar 3
9152 byarna 3
9153 bygga 64
9154 byggande 3
9155 byggandet 6
9156 byggas 12
9157 byggd 1
9158 byggde 3
9159 byggdes 2
9160 bygge 2
9161 bygger 23
9162 bygget 5
9163 byggets 2
9164 bygglåda 1
9165 byggmästare 1
9166 byggnad 10
9167 byggnaden 8
9168 byggnadstillstånd 1
9169 byggnadstillståndet 1
9170 byggs 6
9171 byggstenarna 1
9172 byggt 10
9173 byggts 3
9174 bylte 1
9175 byn 4
9176 byrå 3
9177 byråer 6
9178 byråerna 1
9179 byråkrater 1
9180 byråkraternas 1
9181 byråkrati 22
9182 byråkratin 4
9183 byråkratisk 5
9184 byråkratiska 11
9185 byråkratiskt 4
9186 byrån 5
9187 byråns 1
9188 byta 9
9189 byte 2
9190 byten 1
9191 byter 2
9192 byteshandel 1
9193 bytet 1
9194 bytts 1
9195 byxfickorna 1
9196 byxor 1
9197 byxorna 1
9198 bädd 1
9199 bägare 1
9200 bägge 5
9201 bälte 1
9202 bände 1
9203 bänk 1
9204 bär 36
9205 bära 19
9206 bärande 3
9207 bärare 2
9208 bäras 5
9209 bärighet 1
9210 bärkraft 1
9211 bärs 3
9212 bäst 28
9213 bästa 124
9214 bäste 5
9215 bättra 1
9216 bättre 262
9217 båda 107
9218 bådadera 1
9219 både 186
9220 bågnat 1
9221 bålen 1
9222 bålrullningar 1
9223 bården 1
9224 bås 1
9225 båt 3
9226 båtar 16
9227 båtarna 1
9228 båtarnas 1
9229 båtars 1
9230 båten 1
9231 båtens 2
9232 bébé 1
9233 böcker 11
9234 böckerna 1
9235 böckling 2
9236 böcklingar 2
9237 bödelsdräng 1
9238 böja 1
9239 böjd 1
9240 böjda 1
9241 böjde 5
9242 böjelse 1
9243 böjt 1
9244 bölande 1
9245 bön 1
9246 bönbok 1
9247 bönder 3
9248 bönderna 2
9249 bönen 1
9250 bönens 1
9251 bör 610
9252 börda 4
9253 bördan 7
9254 bördor 1
9255 bördorna 3
9256 börja 123
9257 började 54
9258 början 80
9259 börjar 58
9260 börjat 36
9261 börsen 2
9262 börser 1
9263 börsindex 1
9264 börsmarknaderna 1
9265 börsnoterade 1
9266 börsvärde 2
9267 bössan 1
9268 böter 5
9269 bötesstraff 2
9270 c 2
9271 c'est 1
9272 ca 6
9273 calendas 1
9274 calvinistiska 1
9275 can 1
9276 canapéer 1
9277 canapérecept 1
9278 cancer 2
9279 cancerböld 1
9280 cancerframkallande 1
9281 cannabisen 1
9282 capita 14
9283 case 1
9284 caulerpa 1
9285 cell 2
9286 celler 1
9287 celsius 1
9288 cementerar 2
9289 censurera 1
9290 cent 1
9291 centimeter 3
9292 centra 3
9293 central 29
9294 central- 3
9295 centrala 37
9296 centralafrikanska 1
9297 centralatlanten 1
9298 centralbanken 11
9299 centralbankens 4
9300 centralbanker 1
9301 centralbankerna 1
9302 centraleuropeiska 2
9303 centralförvaltningars 1
9304 centralförvaltningen 1
9305 centralisera 1
9306 centraliserad 2
9307 centraliserade 1
9308 centraliserande 1
9309 centraliserar 2
9310 centraliserat 2
9311 centraliserats 1
9312 centralisering 6
9313 centralistiska 1
9314 centralistiskt 2
9315 centralregering 2
9316 centralregeringen 2
9317 centralstyrningen 1
9318 centralt 10
9319 centre 1
9320 centrerats 1
9321 centrum 27
9322 centrumen 3
9323 ceremonier 1
9324 ceremonin 2
9325 certifiering 1
9326 certifieringssällskap 1
9327 certifikat 3
9328 champagne 2
9329 champagneflaska 1
9330 change 1
9331 chans 30
9332 chansen 7
9333 chanser 5
9334 chanserna 2
9335 chapeau 1
9336 charaderna 1
9337 charmanta 1
9338 charmen 1
9339 chartrar 1
9340 chassid 2
9341 chassiden 3
9342 chassider 2
9343 chassiderna 3
9344 chassidim 1
9345 chassidisk 1
9346 chaufförer 3
9347 check 1
9348 chef 8
9349 chefen 3
9350 chefer 5
9351 cheferna 6
9352 chefs- 1
9353 chefsjobb 1
9354 chefstjänster 1
9355 chilenska 1
9356 chock 1
9357 chockad 2
9358 chocken 3
9359 chocker 1
9360 chockerad 1
9361 chockerade 2
9362 chockerande 4
9363 chockerar 1
9364 chockerna 1
9365 choklad 4
9366 chokladdirektivet 1
9367 chokladvaror 1
9368 cigarett 4
9369 cigaretten 1
9370 cigaretter 2
9371 cigarettmärke 1
9372 cigarettpapper 1
9373 cigarr 1
9374 cigarrask 1
9375 cigarrer 1
9376 cirka 25
9377 cirkel 2
9378 cirkeldiagram 1
9379 cirkelns 1
9380 cirklar 2
9381 cirkulera 1
9382 cirkulerar 5
9383 cirkulerat 1
9384 cirkulärbrev 1
9385 citat 3
9386 citera 10
9387 citerade 1
9388 citerar 20
9389 citeras 3
9390 citrusfrukter 1
9391 civil 7
9392 civil- 1
9393 civila 52
9394 civilbefolkningen 3
9395 civilförsvaret 1
9396 civilförsvarsmakt 1
9397 civilisation 4
9398 civilisationen 1
9399 civilisationens 1
9400 civilisera 1
9401 civiliserad 2
9402 civiliserade 3
9403 civiliserat 4
9404 civilist 1
9405 civilmål 1
9406 civilperson 1
9407 civilpolis 1
9408 civilrätt 1
9409 civilrättens 1
9410 civilrättsligt 1
9411 civilskydd 2
9412 civilskyddet 1
9413 civilt 4
9414 clauses 1
9415 clearingorganisationer 1
9416 close 1
9417 clowneri 1
9418 coccidiostatika 2
9419 cocktailbjudningar 1
9420 cocktailklänning 1
9421 collage 1
9422 cologne 1
9423 combattant 1
9424 comitology 2
9425 commitment 2
9426 common 1
9427 compassion 1
9428 compounder 1
9429 con 1
9430 conditio 2
9431 conduite 1
9432 conference 1
9433 confidence 1
9434 consentiment 1
9435 contradictio 1
9436 contrario 1
9437 contre-filet 1
9438 control 2
9439 copyright 1
9440 corporate 3
9441 corpus 6
9442 correcta 2
9443 correctness 1
9444 cost-benefit-analys 5
9445 costing 1
9446 counter 1
9447 counter-instrument 1
9448 countries 1
9449 coup 1
9450 cowboy 2
9451 creams 1
9452 cricketmatcher 1
9453 crisis 1
9454 cyanid 3
9455 cyanidförgiftat 1
9456 cyanidtillverkning 1
9457 cyberspace 1
9458 cykeln 1
9459 cyklade 1
9460 cyklonen 1
9461 cynisk 1
9462 cynism 1
9463 cyprioter 2
9464 cyprioterna 2
9465 cypriotiska 13
9466 cypriots 1
9467 d 2
9468 d'argent 1
9469 d'essai 1
9470 d'intention 1
9471 da 9
9472 dag 588
9473 dagar 44
9474 dagarna 23
9475 dagarnas 1
9476 dagars 2
9477 dagen 24
9478 dagens 54
9479 daghemsplatser 1
9480 daglig 2
9481 dagliga 15
9482 dagligen 12
9483 dagligt 1
9484 daglönare 1
9485 dagmamma 1
9486 dagordning 42
9487 dagordningen 56
9488 dagordningens 1
9489 dagordnings 1
9490 dagosens 1
9491 dags 39
9492 dagsläget 4
9493 dagstidning 2
9494 dagstidningar 2
9495 dagstidningen 1
9496 dal 1
9497 dalen 2
9498 dalens 2
9499 dam 1
9500 damer 82
9501 damerna 1
9502 damm 8
9503 dammar 5
9504 dammen 2
9505 dammens 1
9506 dammet 1
9507 dammiga 1
9508 dans 3
9509 dansa 2
9510 dansade 1
9511 dansande 1
9512 dansar 2
9513 dansare 1
9514 dansgolvet 1
9515 dansk 5
9516 danska 35
9517 danslektionerna 1
9518 dar 4
9519 darrade 1
9520 dass 1
9521 dasset 1
9522 data 40
9523 databas 3
9524 databasen 3
9525 databasens 1
9526 databaser 5
9527 databasfönstret 3
9528 databasobjekt 2
9529 datablad 8
9530 databladet 2
9531 datadelen 1
9532 dataelement 4
9533 dataexperter 1
9534 datakälla 5
9535 datakällan 3
9536 datamodellen 1
9537 dataområdet 2
9538 dataschemat 1
9539 dataskydd 1
9540 datastrukturen 2
9541 datasäkerhetsrättsligt 1
9542 datatyper 1
9543 datautrustning 1
9544 datavärden 1
9545 dataåtkomstsida 14
9546 dataåtkomstsidan 4
9547 dataåtkomstsidor 3
9548 dataöverföringen 1
9549 daterad 1
9550 dato 1
9551 dator 2
9552 datorbrottslighet 1
9553 datorer 1
9554 datorisering 1
9555 datorn 4
9556 datornät 1
9557 datorskrot 1
9558 datum 21
9559 datumet 4
9560 de 5722
9561 deadline 1
9562 dealt 2
9563 debatt 207
9564 debatten 188
9565 debattens 2
9566 debatter 18
9567 debattera 16
9568 debatterade 4
9569 debatterar 5
9570 debatteras 11
9571 debatterat 4
9572 debatterats 1
9573 debatterna 6
9574 debattinnehållet 2
9575 debattkväll 1
9576 debattskyldigheten 1
9577 debattunderlag 1
9578 debiteras 1
9579 debiterats 1
9580 december 46
9581 december- 1
9582 decemberveckan 1
9583 decennier 9
9584 decennierna 6
9585 decenniers 2
9586 decenniet 5
9587 decennium 7
9588 decentralisera 1
9589 decentraliserad 3
9590 decentraliserade 3
9591 decentraliserar 2
9592 decentraliseras 3
9593 decentraliserat 4
9594 decentralisering 9
9595 decentraliseringen 1
9596 decentraliseringsprocessen 1
9597 decentralistisk 1
9598 definiera 20
9599 definierad 1
9600 definierade 7
9601 definierades 2
9602 definierar 2
9603 definieras 8
9604 definierat 4
9605 definierats 2
9606 definition 23
9607 definitionen 12
9608 definitioner 5
9609 definitionerna 4
9610 definitionsmässigt 5
9611 definitiv 5
9612 definitiva 4
9613 definitivt 17
9614 degenererar 1
9615 degraderas 3
9616 deklaration 1
9617 deklarationen 1
9618 deklarerad 1
9619 deklarerar 1
9620 deklarerats 1
9621 dekor 2
9622 del 385
9623 dela 22
9624 delad 3
9625 delade 9
9626 delades 2
9627 delaktig 3
9628 delaktiga 11
9629 delaktighet 11
9630 delaktigheten 2
9631 delaktigt 2
9632 delar 133
9633 delarna 10
9634 delas 16
9635 delaspekt 1
9636 delat 8
9637 delats 15
9638 delayed 2
9639 delegater 1
9640 delegaterna 2
9641 delegation 22
9642 delegationen 19
9643 delegationens 2
9644 delegationer 4
9645 delegationerna 2
9646 delegations 1
9647 delegera 2
9648 delegeras 3
9649 delegerats 1
9650 delegering 5
9651 delegeringsartikeln 1
9652 delen 77
9653 delfiner 1
9654 delfrågor 1
9655 delgivning 1
9656 delikat 2
9657 dellösning 1
9658 delmängd 1
9659 delmål 1
9660 delning 7
9661 delprivatiseringar 1
9662 delrapporten 1
9663 dels 30
9664 delsession 1
9665 delstater 1
9666 delstaterna 1
9667 delstatsbanker 2
9668 delta 71
9669 deltaga 1
9670 deltagande 74
9671 deltagandet 2
9672 deltagare 4
9673 deltagarinriktade 1
9674 deltagarna 3
9675 deltagarnas 2
9676 deltagit 10
9677 deltar 34
9678 deltid 1
9679 deltidsarbetandets 1
9680 deltidsarbeten 1
9681 deltidssysselsättning 1
9682 deltog 12
9683 delutbetalningen 2
9684 delvis 39
9685 delägarna 1
9686 dem 614
9687 demagoger 1
9688 demagogi 6
9689 demagogiska 1
9690 demaskeras 1
9691 dementera 1
9692 dementerade 1
9693 demilitariseras 1
9694 demilitariseringen 1
9695 demografin 1
9696 demografiska 10
9697 demokrat 5
9698 demokrater 5
9699 demokraterna 1
9700 demokrati 71
9701 demokratier 1
9702 demokratierna 3
9703 demokratiernas 1
9704 demokratifråga 1
9705 demokratin 36
9706 demokratins 8
9707 demokratireform 1
9708 demokratisera 3
9709 demokratisering 3
9710 demokratiseringen 1
9711 demokratiseringens 1
9712 demokratiseringsprocesserna 1
9713 demokratisk 39
9714 demokratiska 102
9715 demokratiskt 40
9716 demoniskt 1
9717 demonstration 7
9718 demonstrationer 4
9719 demonstrationsprojekt 1
9720 demonstrera 3
9721 demonstrerar 1
9722 demonstrerat 1
9723 demontera 2
9724 demontering 3
9725 demonteringen 1
9726 demonteringskraven 1
9727 demonteringsverksamheten 1
9728 den 5944
9729 denied 2
9730 denna 1343
9731 denne 16
9732 dennes 8
9733 densamma 9
9734 densamme 1
9735 departement 3
9736 departementen 5
9737 departementet 2
9738 departementsnivå 1
9739 dependent 1
9740 deponera 1
9741 deponerat 1
9742 deporteringarna 1
9743 depositioner 2
9744 der 9
9745 deras 281
9746 derivat 11
9747 derivaten 2
9748 derivatinstrument 4
9749 derivatives 1
9750 derivatprodukter 1
9751 derivatregleringen 1
9752 des 2
9753 desamma 3
9754 desertering 1
9755 desertörer 1
9756 design 2
9757 designläge 3
9758 designläget 2
9759 designmiljöer 1
9760 designsmiljö 1
9761 desinfektionsmedel 1
9762 desinfektionsmedlet 1
9763 desinficering 1
9764 desperat 6
9765 desperata 3
9766 desperation 1
9767 despoter 1
9768 despotiska 1
9769 dess 268
9770 dessa 941
9771 dessutom 98
9772 dessvärre 9
9773 destabilisera 4
9774 destabiliserande 2
9775 destilleringssamhälle 1
9776 desto 23
9777 destruktiv 2
9778 destruktiva 1
9779 det 9645
9780 detalj 12
9781 detaljanalys 1
9782 detaljbestämmelser 1
9783 detaljdata 3
9784 detaljen 1
9785 detaljer 15
9786 detaljerad 10
9787 detaljerade 16
9788 detaljerat 8
9789 detaljerna 8
9790 detaljflödet 1
9791 detaljfält 1
9792 detaljfälten 1
9793 detaljhandeln 1
9794 detaljkontroll 2
9795 detaljområden 2
9796 detaljområdet 4
9797 detaljplanet 1
9798 detaljproblem 1
9799 detaljreglerade 1
9800 detaljreglering 1
9801 detaljstyr 1
9802 detektiv 1
9803 detektivromaner 1
9804 detektivverksamhet 1
9805 detektorer 1
9806 detonation 1
9807 detsamma 26
9808 detta 2174
9809 det­ 1
9810 devalvering 1
9811 deve 1
9812 development 1
9813 di 1
9814 diagnos 1
9815 diagnosen 1
9816 diagnostik 1
9817 diagram 2
9818 diagrammet 1
9819 diagrammets 1
9820 diagramtyp 1
9821 dialog 66
9822 dialogen 35
9823 dialogens 2
9824 dialoger 1
9825 dialogerna 1
9826 dialogform 1
9827 dialogrutan 1
9828 diamant 1
9829 diamanter 1
9830 diamanterna 2
9831 die 2
9832 diektivförslaget 1
9833 diesel 2
9834 differentierad 3
9835 differentierade 1
9836 differentieras 1
9837 differentierat 1
9838 differentiering 5
9839 differentieringen 2
9840 diffusa 4
9841 différence 1
9842 dig 34
9843 digital 2
9844 digitala 7
9845 diken 1
9846 dikt 1
9847 diktatorer 2
9848 diktatoriska 1
9849 diktatorlärling 1
9850 diktatur 7
9851 diktaturen 2
9852 diktaturer 2
9853 diktaturerna 1
9854 dikter 2
9855 dikterade 1
9856 dikterar 1
9857 dikteras 1
9858 dikterats 1
9859 diktsamlingar 1
9860 dilemma 3
9861 dilemman 1
9862 dilettanteri 1
9863 dill 1
9864 dillkvist 1
9865 dimension 21
9866 dimensionen 16
9867 dimensioner 4
9868 dimensionerna 1
9869 dimma 5
9870 dimman 1
9871 din 6
9872 dina 6
9873 dinehbefolkningen 1
9874 dinehindianerna 4
9875 dinehindianernas 1
9876 dinglade 2
9877 dinglande 1
9878 dioxiderna 1
9879 dioxin 3
9880 dioxinkrisen 2
9881 dioxinskandalen 1
9882 dioxinskräckhistorien 1
9883 dioxinskräckupplevelsen 1
9884 diplomatbeskickningar 1
9885 diplomater 2
9886 diplomati 4
9887 diplomatin 1
9888 diplomatins 1
9889 diplomatisk 5
9890 diplomatiska 12
9891 diplomatiskt 3
9892 diplomatkår 1
9893 direct 1
9894 direkt 112
9895 direkta 17
9896 direktbeskattning 1
9897 direktdialog 2
9898 direktfinansiera 1
9899 direkthjälpen 1
9900 direktinvesteringar 1
9901 direktiv 244
9902 direktiven 16
9903 direktivens 1
9904 direktivet 172
9905 direktivets 16
9906 direktivförslag 2
9907 direktivförslaget 4
9908 direktivtext 1
9909 direktkontakt 1
9910 direktkontakten 1
9911 direktorat 3
9912 direktreaktion 1
9913 direktreklam 3
9914 direktsändes 1
9915 direktsänds 1
9916 direktör 2
9917 direktören 4
9918 direktörens 1
9919 direktörerna 1
9920 direktörstyper 1
9921 dirigera 1
9922 dirigism 1
9923 dis 1
9924 disciplin 9
9925 disciplinerade 1
9926 disciplinering 2
9927 disciplinerna 1
9928 disciplinfrågor 1
9929 disciplinråden 1
9930 disciplinära 4
9931 diset 1
9932 disk 1
9933 diska 1
9934 diskbänken 1
9935 disken 5
9936 diskho 1
9937 diskret 3
9938 diskreta 1
9939 diskretion 1
9940 diskriminera 1
9941 diskriminerade 3
9942 diskriminerande 4
9943 diskrimineras 1
9944 diskriminering 59
9945 diskrimineringar 2
9946 diskrimineringen 3
9947 diskrimineringsförslag 1
9948 diskrimineringskategori 1
9949 diskrimineringskategorierna 1
9950 diskursen 1
9951 diskussion 47
9952 diskussionen 36
9953 diskussioner 47
9954 diskussionerna 13
9955 diskussions- 1
9956 diskussionsdokument 1
9957 diskussionsforum 1
9958 diskussionsgrupp 1
9959 diskussionsprocess 1
9960 diskussionspunkt 1
9961 diskussionspunkten 1
9962 diskussionsunderlag 2
9963 diskussionsämne 2
9964 diskussionsämnen 1
9965 diskutabelt 2
9966 diskutabla 2
9967 diskutera 77
9968 diskuterade 16
9969 diskuterades 4
9970 diskuterar 64
9971 diskuteras 25
9972 diskuterat 19
9973 diskuterats 10
9974 dispenser 1
9975 disponerar 1
9976 disponeras 1
9977 disponibla 2
9978 dispositioner 1
9979 dispositionerna 2
9980 disproportion 1
9981 dispyt 1
9982 disrupters 1
9983 distans 2
9984 distansförhöret 1
9985 distanshandel 1
9986 distinktion 3
9987 distraheras 1
9988 distraktion 1
9989 distribuera 1
9990 distribuerar 2
9991 distribution 3
9992 distributionen 1
9993 distributionsnätens 1
9994 distributionssektorn 1
9995 distributörers 1
9996 distriktsdomare 1
9997 distriktskommissarien 2
9998 dit 38
9999 dithän 1
10000 dithörande 1
10001 ditt 3
10002 ditupp 1
10003 divaner 1
10004 diverse 14
10005 diversehandeln 1
10006 diversifiera 1
10007 diversifierade 1
10008 diversifierat 1
10009 diversifiering 1
10010 divisioner 1
10011 djungel 2
10012 djungeln 1
10013 djungelns 2
10014 djup 11
10015 djupa 12
10016 djupare 8
10017 djupaste 3
10018 djupet 10
10019 djupgående 13
10020 djuphavsfiske 1
10021 djupnade 3
10022 djupnande 1
10023 djupsinnighet 2
10024 djupt 26
10025 djur 14
10026 djur- 5
10027 djurarter 2
10028 djuren 3
10029 djurens 5
10030 djuret 2
10031 djurfoder 25
10032 djurfoderblandningar 1
10033 djurfoderbranschen 1
10034 djurfoderindustrins 1
10035 djurfoderproducenterna 1
10036 djurfodret 3
10037 djurhälsovillkor 1
10038 djurhållningen 1
10039 djurliv 2
10040 djurlivet 1
10041 djurläkemedel 1
10042 djurs 2
10043 djärv 3
10044 djärva 5
10045 djärvare 2
10046 djärvhet 2
10047 djärvt 2
10048 djävlar 1
10049 djävlarna 1
10050 djävul 4
10051 djävulen 1
10052 djävulens 1
10053 djävulska 1
10054 dock 267
10055 dockor 2
10056 doft 3
10057 doftande 1
10058 doften 1
10059 dog 11
10060 dogm 1
10061 dogmatiska 1
10062 dogmen 1
10063 doktor 1
10064 doktrin 4
10065 doktrinen 1
10066 dokument 98
10067 dokumentation 1
10068 dokumentationen 1
10069 dokumenten 8
10070 dokumenterade 1
10071 dokumentet 18
10072 dokumentets 1
10073 dokumentkategorier 1
10074 dokumentskåp 1
10075 dold 3
10076 dolda 1
10077 dollar 18
10078 dollarn 3
10079 dollartecken 1
10080 dolomiten 1
10081 dolt 2
10082 dom 20
10083 domar 8
10084 domare 11
10085 domaren 2
10086 domarkollegier 1
10087 domarna 7
10088 domarnas 1
10089 domen 3
10090 dominans 3
10091 dominansen 1
10092 dominera 3
10093 dominerades 1
10094 dominerande 12
10095 dominerar 1
10096 domineras 4
10097 domino 1
10098 dominospel 1
10099 domkretsar 1
10100 domslut 3
10101 domsrätt 1
10102 domsrätten 1
10103 domstol 13
10104 domstolar 14
10105 domstolarna 11
10106 domstolars 2
10107 domstolen 24
10108 domstolens 7
10109 domstolsavgörande 1
10110 domstolsfall 1
10111 domstolsförhandlingar 2
10112 domstolsförhandlingarna 1
10113 domstolskandidat 1
10114 domstolsmyndighet 1
10115 domstolsprocessen 1
10116 domstolssystemet 2
10117 domstolstvister 1
10118 domstolsutslag 1
10119 domstolsväsen 1
10120 domäner 1
10121 donator 1
10122 donne 1
10123 donor 1
10124 doppade 1
10125 dos 1
10126 dosis 1
10127 dossier 1
10128 dossieren 1
10129 dot.com-företag 1
10130 dotter 3
10131 dotterdirektiv 1
10132 dov 1
10133 dra 75
10134 drabba 3
10135 drabbade 44
10136 drabbades 9
10137 drabbar 13
10138 drabbas 20
10139 drabbat 11
10140 drabbats 21
10141 drack 4
10142 drag 9
10143 dragande 2
10144 dragbilen 1
10145 dragen 6
10146 draget 2
10147 draggade 1
10148 dragit 8
10149 dragits 4
10150 dragna 1
10151 dragningskraft 1
10152 dragspel 1
10153 drake 1
10154 drakgödsel 1
10155 drakonisk 1
10156 dramat 1
10157 dramatiken 1
10158 dramatiserar 1
10159 dramatisk 6
10160 dramatiska 13
10161 dramatiskt 8
10162 draperi 1
10163 draperiet 1
10164 drar 34
10165 dras 6
10166 drastisk 2
10167 drastiska 4
10168 drastiskt 8
10169 dravel 1
10170 drev 7
10171 drevs 3
10172 dricka 7
10173 drickande 1
10174 drickas 1
10175 drickat 1
10176 dricker 4
10177 dricks 1
10178 dricks- 1
10179 dricksvatten 10
10180 dricksvattenförsörjning 1
10181 dricksvattenförsörjningen 2
10182 dricksvattenkvalitet 1
10183 dricksvattnet 2
10184 drift 4
10185 driften 1
10186 driftiga 1
10187 driftighet 1
10188 driftsförhållanden 1
10189 driftsverksamhet 1
10190 driftsvillkoren 1
10191 driftsäkerhet 1
10192 drink 3
10193 drinken 1
10194 driva 29
10195 drivande 3
10196 drivas 2
10197 driver 16
10198 drivfjäder 1
10199 drivfjädern 1
10200 drivgarn 3
10201 driving 1
10202 drivit 2
10203 drivkraft 6
10204 drivkraften 1
10205 drivkrafter 2
10206 drivkrafterna 1
10207 drivmotor 1
10208 drivs 6
10209 drog 26
10210 drogberoende 4
10211 drogeffekter 1
10212 droger 1
10213 drogkulturen 1
10214 drogs 5
10215 droit 2
10216 droppade 1
10217 droppe 3
10218 droppen 2
10219 drottning 2
10220 drottningens 1
10221 drottninglik 1
10222 druckit 3
10223 drucknes 1
10224 drunkna 2
10225 drunknade 2
10226 drunknar 1
10227 drunknat 2
10228 dryck 1
10229 drycker 5
10230 dryckerna 1
10231 dryfta 2
10232 dryftar 2
10233 drygt 8
10234 drägligare 1
10235 drägligt 1
10236 drämde 1
10237 dränka 1
10238 dränkte 2
10239 dråpslag 1
10240 dröja 4
10241 dröjde 3
10242 dröjer 5
10243 dröjsmål 6
10244 dröjt 2
10245 dröm 1
10246 drömde 2
10247 drömma 3
10248 drömmande 1
10249 drömmar 3
10250 drömmen 4
10251 drömtillfälle 1
10252 du 220
10253 dualiseras 1
10254 dubbel 5
10255 dubbelbeskattning 1
10256 dubbeldörrarna 1
10257 dubbelfinansiering 1
10258 dubbelhaka 1
10259 dubbelkontrollera 1
10260 dubbelmoral 1
10261 dubbelrunda 1
10262 dubbelskrovet 2
10263 dubbelt 4
10264 dubbelväggigt 1
10265 dubbla 21
10266 dubblera 3
10267 dubblerade 1
10268 dubbleringar 1
10269 dubbleringen 1
10270 ducka 1
10271 duga 1
10272 duger 1
10273 dugligheten 1
10274 duk 1
10275 dukade 2
10276 dukar 1
10277 dukat 1
10278 duktig 1
10279 duktiga 2
10280 duktigt 1
10281 dum 4
10282 dumhet 3
10283 dumheter 2
10284 dumpades 1
10285 dumpandet 1
10286 dumpning 9
10287 dumt 5
10288 dunans 1
10289 dunder 1
10290 dungen 1
10291 dungens 1
10292 dunkande 2
10293 dunkel 1
10294 dunkelt 1
10295 dunklet 1
10296 dunmjuka 1
10297 duns 1
10298 dures 1
10299 duschade 1
10300 dussin 2
10301 dvala 1
10302 dvs 3
10303 dvs. 125
10304 dy 1
10305 dygder 1
10306 dygn 1
10307 dygnet 1
10308 dyka 4
10309 dyker 8
10310 dykningen 1
10311 dykt 5
10312 dylika 5
10313 dylikt 1
10314 dynamik 7
10315 dynamiken 1
10316 dynamisk 8
10317 dynamiska 10
10318 dynamiskt 2
10319 dynamitladdning 1
10320 dyngbaggar 1
10321 dynggrepen 1
10322 dyningen 1
10323 dyr 3
10324 dyra 3
10325 dyrare 4
10326 dyraste 2
10327 dyrbar 2
10328 dyrbart 1
10329 dyrka 1
10330 dyrkan 1
10331 dyrt 5
10332 dyster 3
10333 dystert 2
10334 dystra 4
10335 däck 3
10336 däckfabrikant 1
10337 däggdjur 2
10338 dämpa 4
10339 dämpad 1
10340 dämpades 1
10341 dämpar 1
10342 dämpas 1
10343 där 906
10344 därav 7
10345 därefter 27
10346 däremellan 1
10347 däremot 39
10348 därför 507
10349 därhemma 1
10350 därhän 3
10351 däri 1
10352 däribland 15
10353 därifrån 8
10354 därigenom 33
10355 därinne 1
10356 därmed 109
10357 därnere 1
10358 däromkring 1
10359 därpå 6
10360 därtill 3
10361 därutanför 1
10362 därute 3
10363 därvid 5
10364 då 486
10365 dåd 1
10366 dådet 1
10367 dålig 14
10368 dåliga 21
10369 dåligt 20
10370 dån 1
10371 dånade 1
10372 dånande 1
10373 dånet 1
10374 dåvarande 3
10375 défense 2
10376 démocratique 1
10377 dö 7
10378 död 25
10379 döda 27
10380 dödade 10
10381 dödades 2
10382 dödande 1
10383 dödar 6
10384 dödas 6
10385 dödat 2
10386 dödats 3
10387 döde 1
10388 döden 3
10389 dödens 3
10390 dödfödd 1
10391 dödhet 1
10392 dödliga 2
10393 dödlighet 1
10394 dödläge 1
10395 dödsdomen 1
10396 dödsdömd 1
10397 dödsfall 2
10398 dödsfallen 2
10399 dödsfrekvensen 1
10400 dödskallar 1
10401 dödskampen 1
10402 dödsliknande 1
10403 dödsmärkt 1
10404 dödsoffer 1
10405 dödsrikets 1
10406 dödsstraff 4
10407 dödsstraffet 8
10408 döende 1
10409 dög 1
10410 dök 12
10411 dölja 21
10412 döljer 11
10413 döljs 4
10414 döma 19
10415 dömande 1
10416 dömas 2
10417 dömd 1
10418 dömda 2
10419 dömde 2
10420 dömer 2
10421 döms 1
10422 dömts 2
10423 döpa 1
10424 döper 3
10425 döpte 1
10426 dör 13
10427 dörr 9
10428 dörrar 6
10429 dörrarna 3
10430 dörrarnas 1
10431 dörren 32
10432 dörrhandtag 1
10433 dörrklockan 1
10434 dörrvredet 1
10435 dörröppningen 1
10436 dörröverstycken 1
10437 dött 12
10438 döttrar 1
10439 döttrarna 1
10440 döva 3
10441 e 4
10442 e-Europa 3
10443 e-Europe 2
10444 e-företagande 1
10445 e-företagandet 1
10446 e-handel 1
10447 e-handeln 6
10448 e-handelsmöjligheter 1
10449 e-mail 1
10450 e-post 4
10451 e-posthastighet 1
10452 e-sidan 1
10453 e.d. 1
10454 eau 1
10455 ebben 4
10456 ebbremsa 1
10457 ecu 6
10458 ed 1
10459 eden 1
10460 effekt 29
10461 effekten 13
10462 effekter 42
10463 effekterna 30
10464 effektfull 1
10465 effektiv 77
10466 effektiva 43
10467 effektivare 34
10468 effektivaste 3
10469 effektivisera 7
10470 effektivisering 2
10471 effektivitet 33
10472 effektiviteten 17
10473 effektivitetsargument 1
10474 effektivitetskriterier 1
10475 effektivitetssprång 1
10476 effektivt 81
10477 effektstudie 1
10478 effektuera 1
10479 efter 493
10480 efterbilda 1
10481 efterbildar 1
10482 efterblivna 1
10483 efterforskningar 4
10484 efterfrågan 18
10485 efterfrågans 1
10486 efterfrågar 2
10487 efterfrågat 1
10488 efterfrågats 2
10489 efterfråge-elasticitet 2
10490 efterfrågningar 1
10491 efterföljande 4
10492 efterföljare 1
10493 efterföljarna 1
10494 eftergift 1
10495 eftergifter 5
10496 eftergivenhet 4
10497 eftergivenheten 1
10498 eftergivna 1
10499 eftergymnasial 1
10500 efterhand 11
10501 efterhandsgranskning 1
10502 efterhandskontrollen 1
10503 efterkommande 1
10504 efterkälken 3
10505 efterlevas 2
10506 efterlevnad 6
10507 efterlevs 8
10508 efterlevts 2
10509 efterlikna 2
10510 efterlysa 1
10511 efterlyser 3
10512 efterlyses 1
10513 efterlysning 1
10514 efterlyst 1
10515 efterlämnade 1
10516 eftermiddag 17
10517 eftermiddagarna 1
10518 eftermiddagen 5
10519 eftermiddagens 1
10520 eftermiddags 3
10521 eftermiddagskaffe 1
10522 eftermiddan 1
10523 eftermäle 1
10524 efterrättstårta 1
10525 eftersatta 11
10526 eftersatthet 3
10527 eftersatthetskriteriet 1
10528 eftersläpning 4
10529 eftersläpningen 1
10530 eftersom 559
10531 eftersträva 6
10532 eftersträvade 6
10533 eftersträvansvärda 1
10534 eftersträvansvärt 1
10535 eftersträvar 9
10536 eftersträvas 5
10537 eftersträvat 1
10538 eftertanke 7
10539 eftertraktade 1
10540 eftertraktar 1
10541 eftertryck 5
10542 eftertryckligen 5
10543 efterträdare 1
10544 efterträdaren 1
10545 efterträdde 1
10546 eftertänksamhet 1
10547 efterverkningar 1
10548 efteråt 7
10549 egen 108
10550 egenansvar 1
10551 egenart 1
10552 egendom 6
10553 egendomen 1
10554 egendomlig 2
10555 egendomligheter 1
10556 egendomligt 5
10557 egendoms 1
10558 egendomsrätt 1
10559 egenföretagande 1
10560 egenföretagare 3
10561 egenföretagarna 1
10562 egenhet 2
10563 egenintresse 1
10564 egenskap 51
10565 egenskapen 11
10566 egenskaper 7
10567 egenskaperna 2
10568 egenskapsinställningarna 1
10569 egentlig 2
10570 egentliga 5
10571 egentligen 121
10572 egentligt 1
10573 eget 75
10574 egg 1
10575 eggande 1
10576 egna 126
10577 egoism 1
10578 egoistiska 4
10579 egyptiska 3
10580 egyptiskt 1
10581 ej 40
10582 ekade 1
10583 ekologisk 8
10584 ekologiska 27
10585 ekologiskt 10
10586 ekon 1
10587 ekonom 1
10588 ekonomer 1
10589 ekonomernas 1
10590 ekonometriska 1
10591 ekonomi 92
10592 ekonomi- 2
10593 ekonomier 17
10594 ekonomierna 7
10595 ekonomiernas 1
10596 ekonomin 74
10597 ekonomins 9
10598 ekonomisk 151
10599 ekonomiska 397
10600 ekonomiske 1
10601 ekonomiskt 83
10602 ekonomiskt-finansiellt 1
10603 ekonomistyrning 9
10604 ekonomistyrningen 4
10605 ekonomisystemet 1
10606 ekosocial 1
10607 ekosystem 8
10608 ekosystemen 6
10609 ekosystemet 5
10610 ekoturism 1
10611 ekvation 1
10612 ekvatorn 1
10613 ekvilibristik 1
10614 el 1
10615 el- 3
10616 el-Sheikh 3
10617 el-Sheikh-avtalet 1
10618 elak 1
10619 elasticitet 1
10620 eld 2
10621 eldade 1
10622 elden 6
10623 eldkvast 1
10624 eldsken 1
10625 eldskenet 2
10626 eldslåga 1
10627 eldstaden 1
10628 eldsvådan 1
10629 electronic 1
10630 elefant 1
10631 elegant 1
10632 elektricitet 3
10633 elektriskt 6
10634 elektrochock 1
10635 elektronik- 1
10636 elektronikavfall 1
10637 elektronikbranschen 1
10638 elektronikindustrin 1
10639 elektronisk 8
10640 elektroniska 13
10641 elektroniskt 9
10642 element 23
10643 elementet 3
10644 elementnamn 1
10645 elementära 5
10646 elevhemmets 1
10647 elfenben 2
10648 elfte 2
10649 eliminera 11
10650 eliminerade 1
10651 eliminerar 1
10652 elimineras 1
10653 eliminerats 1
10654 eliminering 1
10655 elit 3
10656 eliten 1
10657 elits 1
10658 elitutbildning 1
10659 elkostnaderna 1
10660 elle 1
10661 eller 1216
10662 elmaster 1
10663 eloge 2
10664 elräkningar 1
10665 elva 8
10666 elände 1
10667 eländet 1
10668 eländig 2
10669 eländiga 1
10670 emalj 1
10671 emanciperad 1
10672 embargo 2
10673 embargot 5
10674 emblem 1
10675 emblemet 1
10676 embryo 1
10677 embryoform 1
10678 embryostadiet 1
10679 emedan 1
10680 emellan 14
10681 emellanåt 3
10682 emellertid 167
10683 emigration 1
10684 emigrera 2
10685 emissionsgarantier 1
10686 emot 162
10687 emotionell 1
10688 emotionella 1
10689 emotionellt 2
10690 emotser 1
10691 empiriskt 1
10692 en 8226
10693 en-mängd 1
10694 ena 109
10695 enad 2
10696 enade 16
10697 enades 3
10698 enahanda 1
10699 enande 1
10700 enandet 2
10701 enar 1
10702 enas 9
10703 enastående 9
10704 enat 2
10705 enats 8
10706 enbart 94
10707 encefalopati 1
10708 end 1
10709 enda 183
10710 endast 212
10711 endaste 1
10712 ende 3
10713 endemisk 2
10714 endemiska 1
10715 endocrine 1
10716 endogen 1
10717 endogena 1
10718 ene 2
10719 energi 34
10720 energi- 1
10721 energiagenturer 1
10722 energianvändning 6
10723 energibesparing 3
10724 energibesparingar 1
10725 energicentra 1
10726 energidistribution 1
10727 energieffektiva 1
10728 energieffektivitet 2
10729 energier 2
10730 energierna 1
10731 energiformer 1
10732 energiförbrukningen 1
10733 energiförråden 1
10734 energiförsörjning 1
10735 energiförsörjningen 1
10736 energiförsörjningssystem 1
10737 energiimport 2
10738 energikapacitet 1
10739 energikontrollsystem 1
10740 energikrävande 1
10741 energikälla 2
10742 energikällor 34
10743 energikällorna 4
10744 energikällornas 1
10745 energimarknaden 1
10746 energimixen 1
10747 energin 4
10748 energinäten 2
10749 energiområdet 1
10750 energipolitiken 2
10751 energipotential 1
10752 energiproduktion 2
10753 energiproduktionen 1
10754 energiprogram 1
10755 energiprogrammets 1
10756 energiresurser 1
10757 energisektor 1
10758 energisektorerna 1
10759 energisektorn 4
10760 energisk 1
10761 energiska 1
10762 energiskt 3
10763 energisnåla 1
10764 energiutvinning 1
10765 energiåtervinning 1
10766 energiöverföring 1
10767 enerverande 1
10768 enes 1
10769 enfaldiga 1
10770 enformig 1
10771 enformighet 1
10772 engagemang 43
10773 engagemanget 4
10774 engagera 14
10775 engagerad 2
10776 engagerade 11
10777 engagerar 9
10778 engageras 3
10779 engagerat 4
10780 engelsk 2
10781 engelsk-franska 1
10782 engelska 27
10783 engelskspråkiga 1
10784 engelskt 2
10785 engelsman 2
10786 engelsmannen 1
10787 engelsmän 2
10788 engelsmännen 1
10789 engångsåtgärder 1
10790 enhet 19
10791 enheten 4
10792 enheter 12
10793 enheterna 6
10794 enhetlig 27
10795 enhetliga 15
10796 enhetlighet 8
10797 enhetligt 17
10798 enhetsakten 1
10799 enhetschefer 3
10800 enhetscheferna 1
10801 enhetsorganisationen 2
10802 enhetspolitiska 1
10803 enhetspris 1
10804 enhetsstat 1
10805 enhällig 3
10806 enhälliga 4
10807 enhällighet 20
10808 enhälligheten 2
10809 enhällighetsprincip 1
10810 enhällighetsprincipen 2
10811 enhälligt 27
10812 enig 2
10813 eniga 6
10814 enighet 18
10815 enigheten 1
10816 enigt 1
10817 enkel 17
10818 enkelhet 1
10819 enkelhetens 1
10820 enkelmajoritet 1
10821 enkelriktat 1
10822 enkelt 87
10823 enkelväggigt 2
10824 enkla 21
10825 enklare 8
10826 enklast 1
10827 enklaste 2
10828 enlighet 113
10829 enligt 280
10830 enmansföretag 1
10831 enorm 20
10832 enorma 48
10833 enormt 25
10834 enpartisystemet 1
10835 ens 71
10836 ensam 10
10837 ensamma 14
10838 ensamrätt 2
10839 ensamrätten 1
10840 ensamstående 2
10841 ensamt 4
10842 ense 8
10843 ensidig 4
10844 ensidiga 2
10845 ensidigt 8
10846 enskild 15
10847 enskilda 65
10848 enskildas 2
10849 enskilde 5
10850 enskildhet 1
10851 enskildheter 1
10852 enskilt 13
10853 enstaka 11
10854 entiteten 1
10855 entiteter 1
10856 entreprenad 2
10857 entreprenadföretag 1
10858 entreprenör 1
10859 entreprenören 1
10860 entreprenörerna 2
10861 entreprenörsandan 1
10862 entreprenörskap 3
10863 entreprises 2
10864 enträgen 1
10865 enträget 1
10866 entréhallen 1
10867 entusiasm 11
10868 entusiasmen 1
10869 entusiasmerande 2
10870 entusiastisk 1
10871 entusiastiskt 2
10872 entydig 1
10873 entydiga 3
10874 entydigt 6
10875 envar 1
10876 envetenheten 1
10877 envetet 1
10878 envis 1
10879 envisades 3
10880 envisas 2
10881 envishet 6
10882 envist 4
10883 enväldig 1
10884 enögd 1
10885 epidemier 3
10886 episoden 1
10887 epok 4
10888 epoken 2
10889 epokgörande 1
10890 er 568
10891 era 100
10892 erbjuda 29
10893 erbjudande 1
10894 erbjudanden 2
10895 erbjudandet 1
10896 erbjudas 3
10897 erbjuder 25
10898 erbjudit 1
10899 erbjudits 2
10900 erbjuds 6
10901 erbjöd 6
10902 erbjöds 1
10903 erfara 3
10904 erfaren 1
10905 erfarenhet 28
10906 erfarenheten 4
10907 erfarenheter 40
10908 erfarenheterna 10
10909 erfarenhetsutbyte 5
10910 erfarenhetsutbytet 2
10911 erfarit 2
10912 erfarna 1
10913 erfor 1
10914 erforderlig 3
10915 erforderliga 7
10916 erhalten 1
10917 erhålla 4
10918 erhållande 1
10919 erhåller 3
10920 erhållit 7
10921 erhållits 1
10922 erhöll 4
10923 erinra 28
10924 erinrade 7
10925 erinran 1
10926 erinrar 6
10927 erinras 2
10928 erkänd 8
10929 erkända 4
10930 erkände 6
10931 erkändes 2
10932 erkänds 1
10933 erkänna 29
10934 erkännande 31
10935 erkännandet 5
10936 erkännas 8
10937 erkänner 25
10938 erkänns 5
10939 erkänt 3
10940 erkänts 2
10941 eroderar 1
10942 ersatt 3
10943 ersatta 1
10944 ersatts 3
10945 ersätta 30
10946 ersättas 8
10947 ersätter 6
10948 ersättning 16
10949 ersättningar 4
10950 ersättningarna 1
10951 ersättningen 2
10952 ersättningsansvar 2
10953 ersättningsansvaret 1
10954 ersättningsbeloppet 1
10955 ersättningsmedel 1
10956 ersättningsnivåerna 1
10957 ersättningssystemet 1
10958 ersätts 3
10959 ert 136
10960 erövra 2
10961 erövrades 1
10962 erövrar 1
10963 erövrare 1
10964 erövring 1
10965 erövringen 1
10966 erövringståg 1
10967 es 1
10968 eskorteras 1
10969 esogena 1
10970 esprit 1
10971 essensen 1
10972 essere 1
10973 essäer 1
10974 est 1
10975 esterno 2
10976 estetiska 1
10977 estraden 1
10978 et 3
10979 etablera 9
10980 etablerad 3
10981 etablerade 6
10982 etablerar 2
10983 etablerat 2
10984 etablerats 2
10985 etablering 3
10986 etableringskriteriet 1
10987 etablissemangets 1
10988 etapp 6
10989 etappen 3
10990 etapper 4
10991 etappvis 1
10992 etc 1
10993 etc. 11
10994 etik 1
10995 etikett 3
10996 etiketten 1
10997 etisk 1
10998 etiska 2
10999 etiskt 1
11000 etnisk 11
11001 etniska 27
11002 etniskt 8
11003 ett 4558
11004 etthundranio 1
11005 ettåriga 1
11006 ettårsplanen 1
11007 euro 123
11008 euro-staterna 1
11009 euro-äventyret 1
11010 eurofederalistiska 2
11011 euron 42
11012 eurons 6
11013 euroområdet 4
11014 europaparlamentariker 2
11015 europapatent 1
11016 europatjänsteman 1
11017 europavänlig 1
11018 europeiseras 1
11019 europeisering 1
11020 europeisk 222
11021 europeiska 576
11022 europeiske 4
11023 europeiskt 60
11024 europeistisk 1
11025 europrojektet 1
11026 europé 6
11027 européen 1
11028 européer 27
11029 européerna 8
11030 européernas 3
11031 européers 2
11032 euror 2
11033 eurosedlar 1
11034 euroskeptikerna 1
11035 euroskeptiska 1
11036 eurosymboler 1
11037 eutrofiering 1
11038 evakueras 1
11039 evalueringsbefogenheter 1
11040 evenemang 2
11041 eventuell 16
11042 eventuella 32
11043 eventuellt 38
11044 evig 1
11045 eviga 3
11046 evighet 2
11047 evigt 4
11048 ex 10
11049 exakt 44
11050 exakta 17
11051 exakthet 3
11052 examen 5
11053 examensbevis 1
11054 examensbevisen 1
11055 examination 1
11056 examineringsformer 1
11057 examineringskraven 5
11058 examineringsorganen 1
11059 examineringsorganet 1
11060 examineringsvillkoren 1
11061 excellence 1
11062 exceptionell 3
11063 exceptionellt 5
11064 exempel 293
11065 exempelvis 81
11066 exemplar 7
11067 exemplarisk 1
11068 exemplariska 1
11069 exemplariskt 3
11070 exemplen 6
11071 exemplet 11
11072 exigé 1
11073 exilregeringen 1
11074 exiltibetanerna 1
11075 existens 6
11076 existensberättigande 1
11077 existensen 1
11078 existenser 2
11079 existensrätten 1
11080 existentiella 1
11081 existera 7
11082 existerade 1
11083 existerande 6
11084 existerar 27
11085 exklusiv 2
11086 exklusiva 5
11087 exklusivt 1
11088 exkrementer 1
11089 exotiska 1
11090 expandera 4
11091 expanderande 1
11092 expanderar 2
11093 expansion 1
11094 expansionistiska 1
11095 expansionspolitik 1
11096 expansiva 1
11097 expeditionskommission 1
11098 experiment 3
11099 experimentella 1
11100 experimentera 1
11101 experimentet 1
11102 experimentroll 1
11103 experimentstadiet 2
11104 expert 1
11105 experten 1
11106 experter 15
11107 experterna 10
11108 expertgrupp 2
11109 expertgruppen 2
11110 expertgruppens 2
11111 experthjälp 1
11112 expertis 3
11113 expertkommitté 4
11114 expertkommittén 12
11115 expertkommitténs 4
11116 expertkunskap 1
11117 expertrapport 1
11118 expertregeringar 1
11119 expertutskott 1
11120 explicit 2
11121 exploatera 1
11122 exploateras 2
11123 exploaterbara 1
11124 exploatering 3
11125 exploateringen 2
11126 explodera 1
11127 exploderade 1
11128 exploderar 2
11129 explosion 3
11130 explosionen 2
11131 explosionsartad 1
11132 explosionsrisk 1
11133 explosiv 1
11134 exponentiell 3
11135 exponerar 1
11136 exponeras 1
11137 export 8
11138 exportbidrag 1
11139 exportbidragssystemet 1
11140 exportbranscherna 1
11141 exporten 8
11142 exportera 13
11143 exporterar 6
11144 exporteras 4
11145 exporterat 1
11146 exporterna 1
11147 exportindustrier 1
11148 exportintäkterna 2
11149 exportkrediter 1
11150 exportkreditgarantier 1
11151 exportkreditlicens 1
11152 exportkvot 1
11153 exportör 1
11154 exportörer 2
11155 exportörerna 1
11156 expressbud 1
11157 expressfart 1
11158 expresstjänstesektorn 1
11159 extern 3
11160 externa 19
11161 externt 4
11162 extra 34
11163 extraordinär 1
11164 extraordinära 2
11165 extraordinärt 2
11166 extrarum 1
11167 extrem 1
11168 extrema 7
11169 extremhögern 10
11170 extremhögerns 6
11171 extremism 2
11172 extremistaktioner 1
11173 extremister 2
11174 extremistiska 3
11175 extremistiskt 2
11176 extremsituationer 1
11177 extremt 16
11178 f 1
11179 f.d. 20
11180 fabrik 6
11181 fabriken 6
11182 fabrikens 1
11183 fabriker 5
11184 fabrikerna 1
11185 faciliteter 1
11186 facility 1
11187 facken 1
11188 fackförbund 1
11189 fackföreningar 5
11190 fackföreningarna 4
11191 fackföreningen 1
11192 fackföreningsrörelsen 1
11193 fackföreningsrörelsens 1
11194 fackkunskaper 1
11195 facklan 1
11196 fackliga 3
11197 fackmässig 1
11198 fackrörelsen 1
11199 facktermer 1
11200 fact 1
11201 facto 2
11202 fadder 1
11203 fadern 1
11204 faders 1
11205 failures 1
11206 faire 1
11207 fakta 13
11208 faktabas 1
11209 faktainsamlingsresa 2
11210 faktaunderlag 1
11211 faktisk 3
11212 faktiska 14
11213 faktiskt 142
11214 faktor 25
11215 faktorer 30
11216 faktorerna 2
11217 faktorn 5
11218 faktum 150
11219 faktumet 1
11220 falerner 1
11221 fall 282
11222 falla 7
11223 fallen 11
11224 fallenhet 1
11225 faller 24
11226 fallerar 1
11227 fallet 108
11228 fallfärdiga 1
11229 fallfärdigt 1
11230 fallit 10
11231 fallna 1
11232 fallstudie 1
11233 falsk 4
11234 falska 12
11235 falskheten 1
11236 falskmyntare 1
11237 falskmyntarna 1
11238 falskmynteri 1
11239 falskmyntning 3
11240 falskt 2
11241 familj 9
11242 familje- 2
11243 familjeansvaret 3
11244 familjeenheten 1
11245 familjefader 1
11246 familjeförhållandena 1
11247 familjeförändringar 1
11248 familjejordbruk 3
11249 familjejordbruken 1
11250 familjeliv 1
11251 familjelivet 1
11252 familjemedlem 1
11253 familjen 18
11254 familjens 1
11255 familjeovänliga 1
11256 familjepolitik 2
11257 familjer 25
11258 familjerna 1
11259 familjernas 1
11260 familjeägodelar 1
11261 familjeåterförening 2
11262 famn 2
11263 famnen 2
11264 fanan 1
11265 fanatiska 1
11266 fann 9
11267 fanns 96
11268 fanstyg 1
11269 fantasi 3
11270 fantasibilder 1
11271 fantasier 1
11272 fantasifulla 2
11273 fantasilösa 1
11274 fantasin 3
11275 fantasirik 1
11276 fantastisk 3
11277 fantastiska 10
11278 fantastiskt 7
11279 far 38
11280 fara 27
11281 faran 5
11282 farbar 1
11283 farbror 1
11284 farfarsfars 1
11285 farföräldrar 2
11286 farföräldrars 1
11287 farhågor 10
11288 farkost 2
11289 farkosten 1
11290 farleden 1
11291 farlig 12
11292 farliga 39
11293 farligare 1
11294 farligaste 1
11295 farligheterna 1
11296 farligt 53
11297 farmakologiska 1
11298 farmor 24
11299 farmors 3
11300 farofyllda 1
11301 faror 5
11302 farorna 1
11303 farozon 1
11304 fars 6
11305 farsartade 1
11306 farsot 1
11307 farsoten 1
11308 farsoter 1
11309 fart 8
11310 farten 1
11311 fartyg 61
11312 fartygen 23
11313 fartygens 8
11314 fartyget 16
11315 fartygets 3
11316 fartygs 3
11317 fartygsavfall 1
11318 fartygsbesättningar 1
11319 fartygsgenererade 1
11320 fartygsgenererat 4
11321 fartygsinspektionen 1
11322 fartygsinspektionsbolaget 1
11323 fartygsolyckan 2
11324 fartygsolyckor 1
11325 fartygssidorna 1
11326 fartygsskrov 9
11327 fartygssäkerhet 2
11328 fartygssäkerheten 1
11329 fartygstankrarna 1
11330 fartygsägaren 1
11331 farvatten 14
11332 fas 15
11333 fasa 1
11334 fasaden 1
11335 fasansfull 1
11336 fasansfulla 1
11337 fasat 1
11338 fascineras 1
11339 fascism 2
11340 fascismen 1
11341 fascismens 1
11342 fascistdiktators 1
11343 fascisterna 2
11344 fascisternas 1
11345 fascistisk 1
11346 fascistiska 1
11347 fascistiskt 2
11348 fasen 4
11349 faser 2
11350 faserna 2
11351 fasor 1
11352 fast 96
11353 fasta 18
11354 fasthet 2
11355 fastigheten 1
11356 fastklamrade 1
11357 fastklängda 1
11358 fastkubikmeter 1
11359 fastlagd 1
11360 fastlagda 1
11361 fastlagt 1
11362 fastlagts 2
11363 fastland 2
11364 fastlandet 5
11365 fastlägga 1
11366 fastläggas 1
11367 fastläggs 1
11368 fastnade 1
11369 fastnar 1
11370 fastnat 2
11371 fastsatt 1
11372 fastslagen 1
11373 fastslaget 1
11374 fastslagit 1
11375 fastslagits 2
11376 fastslagna 1
11377 fastslog 4
11378 fastslogs 2
11379 fastslå 9
11380 fastslår 6
11381 fastslås 14
11382 fastställa 60
11383 fastställande 13
11384 fastställandet 4
11385 fastställas 9
11386 fastställd 4
11387 fastställda 8
11388 fastställde 3
11389 fastställdes 10
11390 fastställer 17
11391 fastställs 19
11392 fastställt 5
11393 fastställts 17
11394 fastän 7
11395 fatala 1
11396 fatalitet 1
11397 fatalt 2
11398 fatet 1
11399 fatt 1
11400 fatta 54
11401 fattade 14
11402 fattades 9
11403 fattar 16
11404 fattas 32
11405 fattat 4
11406 fattats 13
11407 fattig 1
11408 fattiga 40
11409 fattigare 6
11410 fattigaste 19
11411 fattigbasaren 2
11412 fattigdom 36
11413 fattigdomen 30
11414 fattigdomsbekämpning 1
11415 fattigdomsbekämpningen 1
11416 fattigdomsbekämpningens 1
11417 fattigdomsdrabbade 1
11418 fattigdomsfokusering 1
11419 fattigdomsgräns 1
11420 fattigdomsgränsen 1
11421 fattigdomsgränser 2
11422 fattigdomsproblematiken 1
11423 fattigdomsproblemen 1
11424 fattigmat 1
11425 fattigt 1
11426 fattning 1
11427 fauna 2
11428 favelas 1
11429 favoritlektyr 1
11430 favör 1
11431 fax 2
11432 faxa 1
11433 feber 1
11434 febrigt 1
11435 februari 48
11436 federal 6
11437 federala 3
11438 federalism 4
11439 federalist 1
11440 federalister 1
11441 federalisterna 1
11442 federalistisk 3
11443 federalistiska 2
11444 federalt 3
11445 federation 3
11446 federationen 2
11447 federationens 1
11448 federationskärna 1
11449 fee 1
11450 fee-system 1
11451 fee-systemet 2
11452 fel 50
11453 felaktig 9
11454 felaktiga 2
11455 felaktigare 1
11456 felaktighet 1
11457 felaktigheter 2
11458 felaktigt 20
11459 felande 1
11460 felar 1
11461 felberäkning 1
11462 felciterad 1
11463 felet 1
11464 felkvot 1
11465 felringning 1
11466 felräkningen 1
11467 felsyn 1
11468 feltolkat 1
11469 felöversättning 2
11470 fem 96
11471 femdubblats 1
11472 femfaldigat 1
11473 femminuterssändning 1
11474 fempunktsprogram 1
11475 femte 21
11476 femtedel 3
11477 femtedelar 1
11478 femtedelen 1
11479 femti 1
11480 femtielfte 1
11481 femtio 10
11482 femtioelfte 1
11483 femtioelva 1
11484 femtiotal 1
11485 femtioårsperiodens 1
11486 femton 37
11487 femtonhundra 1
11488 femtonhundratalet 1
11489 femåriga 1
11490 femårigt 1
11491 femårsperiod 7
11492 femårsperioden 1
11493 femårsplan 2
11494 femårsplanen 5
11495 femårsplaner 2
11496 femårsprogram 8
11497 femårsprogrammet 3
11498 fenomen 12
11499 fenomenet 4
11500 fernissade 1
11501 fest 5
11502 fester 1
11503 festerna 1
11504 festkvällar 1
11505 festligheterna 3
11506 festligt 1
11507 festregeln 1
11508 feststämning 1
11509 feta 2
11510 fiaskona 1
11511 fiaskot 1
11512 fick 149
11513 ficka 1
11514 fickan 3
11515 fickor 1
11516 fickorna 3
11517 fiducia 1
11518 fiende 5
11519 fiender 5
11520 fiendskap 1
11521 fientlig 1
11522 fientliga 3
11523 fientligheterna 3
11524 fientligt 1
11525 figur 1
11526 fikar 1
11527 fil 3
11528 filantropi 1
11529 filen 6
11530 filer 1
11531 filerna 1
11532 filformat 2
11533 filformatet 1
11534 film 1
11535 filmdukar 1
11536 filmen 1
11537 filmens 1
11538 filmer 1
11539 filmsuccé 1
11540 filoberoende 1
11541 filosof 1
11542 filosofi 9
11543 filosofibok 1
11544 filosofin 2
11545 filosofisk 2
11546 filosofiska 2
11547 filtar 3
11548 filten 1
11549 filter 2
11550 filteraxeln 1
11551 filterfunktioner 1
11552 filterfält 3
11553 filterfältet 1
11554 filterområdet 3
11555 filtrera 11
11556 filtrerade 1
11557 filtrerar 4
11558 filtreras 2
11559 filtrerat 2
11560 filtrering 2
11561 filtreringen 1
11562 fin 1
11563 fina 8
11564 finans 1
11565 finans- 1
11566 finansdepartementet 1
11567 finanser 5
11568 finanseringsreformen 1
11569 finanserna 2
11570 finansernas 1
11571 finansföretagens 1
11572 finansgrupp 1
11573 finansiell 12
11574 finansiella 75
11575 finansiellt 17
11576 finansiera 31
11577 finansierad 2
11578 finansierade 3
11579 finansierar 5
11580 finansieras 25
11581 finansierat 2
11582 finansierats 3
11583 finansiering 34
11584 finansieringen 31
11585 finansieringsbeloppet 1
11586 finansieringsbidrag 1
11587 finansieringsinstrument 1
11588 finansieringsinstrumentet 2
11589 finansieringskapital 1
11590 finansieringskällor 1
11591 finansieringsmarknaden 1
11592 finansieringsmetoder 1
11593 finansieringsmodell 1
11594 finansieringsmöjligheter 1
11595 finansieringspaketet 1
11596 finansieringsplan 1
11597 finansieringsplanerna 1
11598 finansieringsprogram 1
11599 finansieringsramar 1
11600 finansieringsramen 1
11601 finansieringsstöd 1
11602 finansieringssystemen 1
11603 finansieringstjänster 1
11604 finansieringsvolym 2
11605 finansieringsåtgärder 1
11606 finansinstituten 2
11607 finansinstrument 1
11608 finansiärer 2
11609 finansiärerna 2
11610 finansmarknaderna 1
11611 finansmarknadernas 1
11612 finansmedlen 1
11613 finansminister 2
11614 finansministern 3
11615 finansministerns 1
11616 finansministrarna 1
11617 finansmän 1
11618 finanspolitik 1
11619 finansprogram 1
11620 finansprotokoll 1
11621 finansprotokollen 2
11622 finansredskap 1
11623 finanssystem 1
11624 finanstekniska 1
11625 finansutskott 1
11626 finaste 2
11627 finding 1
11628 finesse 1
11629 finesser 1
11630 finfördela 1
11631 finge 1
11632 fingeravtrycken 1
11633 fingervisning 2
11634 fingrar 2
11635 fingrarna 4
11636 fingret 2
11637 finhet 1
11638 finkänsliga 1
11639 finkänsligt 1
11640 finländare 1
11641 finländska 9
11642 finna 56
11643 finnas 112
11644 finner 27
11645 finnig 1
11646 finns 924
11647 finsk 4
11648 finska 10
11649 finskuren 1
11650 finskurna 1
11651 fint 2
11652 fira 4
11653 firade 1
11654 firma 1
11655 firman 2
11656 fisk 24
11657 fiska 12
11658 fiskades 1
11659 fiskar 11
11660 fiskare 12
11661 fiskaren 2
11662 fiskarna 10
11663 fiskarnas 2
11664 fiskarter 5
11665 fiskas 1
11666 fiskats 1
11667 fiskbankar 1
11668 fiskbestånd 5
11669 fiskbestånden 5
11670 fiskbeståndet 2
11671 fiske 36
11672 fiske- 3
11673 fiskeansträngningar 1
11674 fiskeansträngningarna 1
11675 fiskeansträngningen 1
11676 fiskeavtalen 1
11677 fiskebankarna 1
11678 fiskebåtar 1
11679 fiskedagarna 1
11680 fiskefartyg 3
11681 fiskefartyget 1
11682 fiskeflotta 2
11683 fiskeflottan 1
11684 fiskeflottor 1
11685 fiskefrågan 1
11686 fiskeindustrins 1
11687 fiskekvoterna 1
11688 fiskelivet 1
11689 fiskemetodernas 1
11690 fiskemängden 1
11691 fiskemöjligheter 4
11692 fisken 8
11693 fiskens 1
11694 fiskeodlingar 1
11695 fiskeområde 1
11696 fiskeområdet 1
11697 fiskeorganisationerna 1
11698 fiskepolitik 1
11699 fiskeprodukter 1
11700 fiskeprodukterna 1
11701 fiskeproduktionen 2
11702 fiskeredskap 2
11703 fiskeredskapen 2
11704 fiskeregion 1
11705 fiskeresurser 1
11706 fiskeresurserna 10
11707 fiskeriansträngningarna 1
11708 fiskeriet 3
11709 fiskerifrågor 1
11710 fiskeriförvaltning 3
11711 fiskeriindustri 1
11712 fiskeriindustrin 1
11713 fiskerikommittén 1
11714 fiskerilagstiftningen 1
11715 fiskerinäring 1
11716 fiskerinäringen 9
11717 fiskerinäringens 1
11718 fiskeriområdet 3
11719 fiskeriorganisation 1
11720 fiskeriorganisationerna 4
11721 fiskeripolitik 10
11722 fiskeripolitiken 35
11723 fiskeripolitikens 2
11724 fiskeriresurserna 1
11725 fiskerisektor 3
11726 fiskerisektorer 1
11727 fiskerisektorn 23
11728 fiskeristatistiken 1
11729 fiskeriutskott 3
11730 fiskeriutskottet 26
11731 fiskeriutskottets 2
11732 fiskeriverksamhet 6
11733 fiskeriverksamheten 6
11734 fiskerättigheter 2
11735 fiskesamhällen 3
11736 fiskesamhällenas 1
11737 fiskesektorer 1
11738 fiskesektorn 4
11739 fiskestopp 1
11740 fisket 39
11741 fisketrycket 3
11742 fiskets 3
11743 fiskeuppgifter 1
11744 fiskevattnen 2
11745 fiskeverksamheten 1
11746 fiskfångst 1
11747 fiskfångstfartyg 1
11748 fiskgrossister 1
11749 fiskodling 3
11750 fiskodlingar 1
11751 fiskodlingen 1
11752 fiskodlingssektorn 1
11753 fiskprodukter 1
11754 fisksjukdomar 2
11755 fission 1
11756 fixa 1
11757 fixera 1
11758 fjol 6
11759 fjolårets 1
11760 fjorton 17
11761 fjortonde 1
11762 fjortonsidiga 1
11763 fjärde 32
11764 fjärde- 1
11765 fjärdedel 2
11766 fjärdedelar 3
11767 fjärilarna 1
11768 fjärma 1
11769 fjärmade 1
11770 fjärran 2
11771 flacka 1
11772 fladdermusliknande 1
11773 fladdrande 2
11774 flagg 10
11775 flagga 4
11776 flaggan 1
11777 flaggens 1
11778 flaggorna 1
11779 flaggskepp 1
11780 flaggstång 1
11781 flagrant 2
11782 flamländska 2
11783 flammade 1
11784 flammat 1
11785 flammorna 1
11786 flampulver 2
11787 flamskyddsmedel 5
11788 flamskyddsmedlen 1
11789 flaska 5
11790 flaskan 3
11791 flaskhals 1
11792 flaskor 2
11793 flaskorna 1
11794 fler 75
11795 flera 217
11796 flerstatlig 1
11797 flertal 12
11798 flertalet 11
11799 flerårig 3
11800 fleråriga 9
11801 flerårigt 8
11802 flerårsbasis 1
11803 flerårsbudget 1
11804 flesta 59
11805 flexibel 14
11806 flexibelt 13
11807 flexibilisering 1
11808 flexibilitet 36
11809 flexibiliteten 3
11810 flexibilitetsklausul 2
11811 flexibla 12
11812 flexiblare 3
11813 flexible 1
11814 flicka 5
11815 flickan 2
11816 flickans 1
11817 flickor 6
11818 flickorna 2
11819 flickors 1
11820 flimret 1
11821 flin 1
11822 flinade 2
11823 flingor 2
11824 flintskallig 1
11825 flirta 1
11826 flit 2
11827 fliten 1
11828 flitigare 1
11829 flock 1
11830 flod 7
11831 flodarm 1
11832 flodbåt 1
11833 floden 27
11834 flodens 1
11835 floder 8
11836 floderna 3
11837 flodernas 2
11838 floders 1
11839 flodledens 1
11840 flodmynningen 3
11841 flodstränder 1
11842 flodstränderna 1
11843 flodvattendistrikt 1
11844 flodvattendistrikten 1
11845 flodvattnet 1
11846 flodvåg 1
11847 flora 2
11848 flottan 5
11849 flottiga 1
11850 flottigt 1
11851 flottkapacitet 1
11852 flottkapaciteten 1
11853 flottorna 2
11854 fluga 1
11855 flugit 1
11856 flugor 1
11857 flutit 1
11858 fly 1
11859 flydde 3
11860 flyg 5
11861 flyga 6
11862 flygande 3
11863 flyganfall 1
11864 flygblad 1
11865 flygbolag 2
11866 flygbombningarna 1
11867 flyger 2
11868 flyget 3
11869 flygkrascherna 1
11870 flyglinjerna 1
11871 flygplan 3
11872 flygplanen 1
11873 flygplanet 1
11874 flygplanskerosin 1
11875 flygplats 2
11876 flygplatsen 3
11877 flygplatser 2
11878 flygpriserna 1
11879 flygräd 1
11880 flygs 1
11881 flygsäkerheten 1
11882 flygtransport 1
11883 flygtransporter 2
11884 flygtransporterna 1
11885 flygturer 1
11886 flygvärdinnan 1
11887 flykt 5
11888 flykten 5
11889 flyktig 1
11890 flykting 2
11891 flykting- 1
11892 flyktingar 30
11893 flyktingarna 8
11894 flyktingeländet 1
11895 flyktingfonden 1
11896 flyktingfrågor 1
11897 flyktingkommissariat 2
11898 flyktingpolitik 3
11899 flyktingpolitiken 2
11900 flyktingstatus 5
11901 flyktingströmmarnas 1
11902 flyktingstödet 1
11903 flyktmöjlighet 1
11904 flyr 1
11905 flyta 1
11906 flytande 1
11907 flyter 2
11908 flytet 1
11909 flytetyg 1
11910 flytt 3
11911 flytta 24
11912 flyttade 7
11913 flyttar 15
11914 flyttas 12
11915 flyttat 5
11916 flyttats 1
11917 flyttfåglar 1
11918 flyttningen 1
11919 flyttningsprogram 1
11920 flyttningsprogrammet 1
11921 fläck 5
11922 fläckar 3
11923 fläcken 2
11924 fläckigt 1
11925 fläkt 1
11926 fläktarna 2
11927 flämtade 3
11928 flämtande 2
11929 fläng 1
11930 flåsande 4
11931 flöde 1
11932 flöden 2
11933 flödet 3
11934 flödiga 1
11935 flög 4
11936 flöjt 1
11937 flörtade 1
11938 flörtig 1
11939 flöt 4
11940 foder 10
11941 foderantibiotika 1
11942 foderblandningar 2
11943 foderdirektivet 1
11944 fodermaterial 1
11945 fodertillsatsen 1
11946 fodertillsatser 14
11947 fodertillsatserna 3
11948 fodertillverkares 1
11949 fog 1
11950 foga 2
11951 fogades 1
11952 fogas 1
11953 fogat 3
11954 foie 3
11955 fokus 5
11956 fokusera 7
11957 fokuserar 7
11958 fokuseras 2
11959 fokuserat 1
11960 fokusering 5
11961 fokuseringen 1
11962 folk 71
11963 folkbibliotek 1
11964 folken 8
11965 folkens 9
11966 folket 27
11967 folketing 1
11968 folketinget 2
11969 folkets 13
11970 folkgrupp 1
11971 folkgrupper 2
11972 folkgrupperna 7
11973 folkhälsa 29
11974 folkhälsan 13
11975 folkhälsans 1
11976 folkhälsoaspekterna 1
11977 folkhälsofråga 2
11978 folkhälsoplanet 1
11979 folkhälsorisk 1
11980 folkhälsoskäl 1
11981 folklagren 2
11982 folklore 1
11983 folkmassan 1
11984 folkmord 7
11985 folkmyllret 2
11986 folkomröstning 5
11987 folkomröstningar 3
11988 folkomröstningen 1
11989 folkopinion 1
11990 folkpartiet 16
11991 folkpartiets 26
11992 folkregeringar 1
11993 folkrepublikens 1
11994 folkräkning 1
11995 folkräkningen 1
11996 folkrätt 1
11997 folkrätten 3
11998 folkrörelserna 1
11999 folks 7
12000 folkskolorna 1
12001 folkstyrets 1
12002 folksägner 1
12003 folktomt 1
12004 folkvalda 12
12005 folkvaldas 1
12006 fond 12
12007 fondandelar 1
12008 fondbolagen 1
12009 fonden 8
12010 fonder 32
12011 fonderna 15
12012 fondernas 1
12013 fondföretag 14
12014 fondföretagen 6
12015 fondföretagens 2
12016 fondföretagsinvesteringar 1
12017 fondförvaltare 2
12018 fondmedel 3
12019 fonduppbyggnad 1
12020 for 15
12021 fora 3
12022 force 3
12023 forcerade 1
12024 fordon 61
12025 fordonen 8
12026 fordonet 2
12027 fordons 1
12028 fordonsindustrin 1
12029 fordonsmärken 1
12030 fordonspark 1
12031 fordonstillverkare 1
12032 fordonstillverkarna 2
12033 fordonsägaren 1
12034 fordonsåtervinningen 1
12035 fordra 1
12036 fordrande 1
12037 fordrar 3
12038 fordras 10
12039 fordringar 1
12040 forell 2
12041 form 102
12042 forma 1
12043 formalism 1
12044 formalitet 2
12045 formaliteter 2
12046 formandet 1
12047 formar 1
12048 format 5
12049 formatering 1
12050 formateringen 3
12051 formationer 1
12052 formatmallar 1
12053 formats 2
12054 formel 3
12055 formell 9
12056 formella 6
12057 formellt 21
12058 formen 7
12059 former 32
12060 formering 1
12061 formerna 6
12062 formulera 10
12063 formulerad 1
12064 formulerade 8
12065 formulerades 2
12066 formuleras 7
12067 formulerat 3
12068 formulerats 6
12069 formulering 7
12070 formuleringar 5
12071 formuleringarna 1
12072 formuleringen 6
12073 formulär 18
12074 formuläret 1
12075 formulärets 2
12076 forna 3
12077 fornminnena 1
12078 forsarna 1
12079 forska 1
12080 forskare 8
12081 forskares 1
12082 forskning 71
12083 forskningen 8
12084 forskningens 2
12085 forsknings- 2
12086 forskningsaktiviteterna 1
12087 forskningsarbeten 1
12088 forskningsbidrag 1
12089 forskningsinformation 1
12090 forskningsinfrastrukturen 1
12091 forskningsområde 4
12092 forskningsområdet 1
12093 forskningsplats 1
12094 forskningspolitik 2
12095 forskningsprogram 5
12096 forskningsprogrammen 1
12097 fort 18
12098 fortare 1
12099 fortbildning 10
12100 fortbildningsprogram 1
12101 fortet 1
12102 fortfarande 296
12103 fortgå 7
12104 fortgående 6
12105 fortlevnad 2
12106 fortlöpande 5
12107 fortlöper 1
12108 fortplantas 1
12109 fortsatt 20
12110 fortsatta 12
12111 fortsatte 16
12112 fortskaffningsmedel 1
12113 fortskrida 1
12114 fortskridande 2
12115 fortskrider 3
12116 fortsätt 2
12117 fortsätta 133
12118 fortsättas 1
12119 fortsätter 76
12120 fortsättning 15
12121 fortsättningen 28
12122 fortsättningsvis 4
12123 forum 8
12124 forumet 5
12125 forêts 1
12126 fosfor 1
12127 fosforrött 1
12128 fossila 2
12129 fosterland 2
12130 fot 5
12131 fotboll 1
12132 fotbollsbedrägerierna 1
12133 fotbollsplan 1
12134 foten 4
12135 fotfäste 1
12136 fotgängarna 1
12137 fotoförstoringar 1
12138 fotograferade 1
12139 fotografi 3
12140 fotografier 2
12141 fotona 1
12142 fots 2
12143 fotspår 2
12144 fotsvamp 1
12145 frack 1
12146 fragment 1
12147 fragmentariskt 1
12148 fragmenterade 1
12149 frakta 1
12150 fraktats 1
12151 fraktens 2
12152 fraktfartyg 1
12153 fraktfordon 1
12154 fram 690
12155 frambesvärja 1
12156 frambringade 1
12157 frambringar 1
12158 framdeles 5
12159 framfart 2
12160 framfusigt 1
12161 framfödde 1
12162 framför 320
12163 framföra 42
12164 framförallt 1
12165 framförande 1
12166 framföranden 3
12167 framföras 1
12168 framförd 1
12169 framförde 13
12170 framförhandlad 1
12171 framförhandlas 1
12172 framförhandlats 1
12173 framförs 7
12174 framfört 12
12175 framförts 17
12176 framgick 4
12177 framgå 3
12178 framgång 44
12179 framgångar 13
12180 framgångarna 2
12181 framgångarnas 1
12182 framgången 7
12183 framgångens 1
12184 framgångsfaktor 1
12185 framgångsrik 19
12186 framgångsrika 12
12187 framgångsrikt 19
12188 framgångssagor 1
12189 framgår 26
12190 framgått 2
12191 framhärda 1
12192 framhärdandet 1
12193 framhärdar 1
12194 framhäva 4
12195 framhävas 2
12196 framhävde 1
12197 framhäver 1
12198 framhävs 1
12199 framhävt 1
12200 framhålla 25
12201 framhållas 2
12202 framhåller 12
12203 framhållit 8
12204 framhålls 2
12205 framhöll 6
12206 framhölls 1
12207 framkalla 2
12208 framkallade 2
12209 framkallar 1
12210 framkallat 5
12211 framkastat 1
12212 framkom 3
12213 framkommer 8
12214 framkommit 7
12215 framlade 1
12216 framlagda 8
12217 framlagt 5
12218 framlagts 6
12219 framlägga 2
12220 framläggandet 3
12221 framlägger 2
12222 framläggs 2
12223 frammana 1
12224 framme 3
12225 framröstade 1
12226 framsida 1
12227 framskjuten 1
12228 framskjutna 2
12229 framskrider 1
12230 framskridet 1
12231 framskridna 1
12232 framsteg 85
12233 framstegen 7
12234 framsteget 2
12235 framstod 1
12236 framställa 9
12237 framställan 1
12238 framställd 1
12239 framställde 1
12240 framställer 1
12241 framställning 10
12242 framställningar 9
12243 framställningarna 1
12244 framställningen 2
12245 framställs 3
12246 framställt 1
12247 framställts 2
12248 framstå 2
12249 framstående 10
12250 framstår 6
12251 framstötar 1
12252 framsätet 2
12253 framtagandet 4
12254 framtagits 1
12255 framtagning 1
12256 framtid 59
12257 framtida 62
12258 framtiden 146
12259 framtidens 4
12260 framtidsbild 1
12261 framtidsdugliga 1
12262 framtidsförmåga 1
12263 framtidshopp 1
12264 framtidsinriktad 1
12265 framtidsinriktat 1
12266 framtidsorienterad 1
12267 framtidsorienterat 1
12268 framtidsutsikter 5
12269 framtidsutsikterna 1
12270 framtoning 1
12271 framträda 2
12272 framträdande 7
12273 framträder 4
12274 framtvingade 1
12275 framtvingar 1
12276 framtvingas 2
12277 framtvingbara 1
12278 framväxande 3
12279 framväxten 1
12280 framåt 66
12281 framåtböjd 1
12282 framåtmarsch 1
12283 framåtskridande 1
12284 framöver 12
12285 franc 5
12286 franca 1
12287 franchisesystem 1
12288 frankiskt 1
12289 fransk 5
12290 franska 75
12291 franske 3
12292 franskt 2
12293 fransktalande 1
12294 franskägt 1
12295 fransmän 1
12296 fransmännen 5
12297 frapperande 1
12298 frasen 1
12299 fraser 1
12300 frasig 1
12301 fred 65
12302 fredag 6
12303 fredagen 3
12304 freden 20
12305 fredens 4
12306 fredlig 13
12307 fredliga 4
12308 fredligt 4
12309 fredsansträngningar 1
12310 fredsavtal 6
12311 fredsavtalen 1
12312 fredsavtalet 4
12313 fredsbeskyddare 1
12314 fredsbevarande 6
12315 fredsbyggande 2
12316 fredsbyggare 1
12317 fredsfrämjande 1
12318 fredsförhandlingarna 3
12319 fredsgrupper 1
12320 fredslösning 1
12321 fredsordning 1
12322 fredsorganisationer 1
12323 fredspartner 1
12324 fredsplan 1
12325 fredsprocess 6
12326 fredsprocessen 37
12327 fredsprocessens 2
12328 fredsprocesser 1
12329 fredsrörelse 1
12330 fredssamarbete 1
12331 fredssamtal 1
12332 fredssamtalen 4
12333 fredssituation 1
12334 fredsskapande 1
12335 fredsstiftande 1
12336 fredsstyrka 1
12337 fredsuppgörelse 3
12338 free 1
12339 frekventera 2
12340 frenetiskt 1
12341 fresker 1
12342 fresta 1
12343 frestas 1
12344 frestelsen 3
12345 fri 47
12346 fri- 32
12347 fria 67
12348 friare 1
12349 friat 1
12350 frid 3
12351 fridfullt 1
12352 fridsamt 1
12353 frigiven 1
12354 frigivningen 1
12355 frigjorda 1
12356 frigjordhet 1
12357 frigjort 1
12358 frigör 1
12359 frigöra 8
12360 frigörande 1
12361 frigöras 1
12362 frigörs 1
12363 frihandel 1
12364 frihandeln 1
12365 frihandelns 4
12366 frihandelsavtalen 1
12367 frihandelsområde 1
12368 frihandelsområden 1
12369 frihandelsområdena 1
12370 frihandelspolitiken 1
12371 frihandelsuppgörelser 1
12372 frihandelsvänliga 1
12373 frihandelszon 1
12374 frihet 97
12375 friheten 20
12376 frihetens 5
12377 friheter 11
12378 friheterna 8
12379 frihetsberövad 1
12380 frihetsberövande 1
12381 frihetskamp 1
12382 frihetskänsla 1
12383 frihetsparti 1
12384 frikostigt 2
12385 friktionsfria 1
12386 frilansande 1
12387 frimärken 1
12388 frimärkspriser 1
12389 frisersalong 1
12390 frisk 2
12391 friska 3
12392 friskt 2
12393 frisläppande 3
12394 frisläppandet 1
12395 frisläppt 1
12396 fristaten 1
12397 fristen 1
12398 frister 2
12399 friställningar 1
12400 fristående 3
12401 fritids- 1
12402 fritidssituationer 1
12403 fritidssysselsättningar 1
12404 fritt 18
12405 frivillig 5
12406 frivillig- 1
12407 frivilliga 14
12408 frivilligas 1
12409 frivilligorganisationer 1
12410 frivilligsektorn 1
12411 frivilligt 7
12412 frodas 6
12413 from 1
12414 fromma 3
12415 front 1
12416 frontalangreppet 1
12417 fronten 4
12418 frontlinjen 1
12419 frosten 1
12420 fru 166
12421 frukost 2
12422 frukostbordet 1
12423 frukosten 2
12424 frukostägg 1
12425 frukt 4
12426 fruktade 3
12427 fruktades 1
12428 fruktan 5
12429 fruktande 1
12430 fruktansvärd 5
12431 fruktansvärda 10
12432 fruktansvärt 5
12433 fruktar 13
12434 fruktat 1
12435 fruktbara 1
12436 fruktbart 7
12437 frukten 2
12438 fruktkaka 1
12439 fruntimmer 1
12440 frusenheten 1
12441 frusna 1
12442 frustade 1
12443 frustar 2
12444 frustration 4
12445 frustrationen 2
12446 frustrerade 1
12447 frustrering 1
12448 frysa 2
12449 fräckhet 1
12450 fräckheten 1
12451 fräkniga 1
12452 fräknigt 1
12453 främja 116
12454 främjade 2
12455 främjande 16
12456 främjandet 11
12457 främjar 32
12458 främjare 1
12459 främjas 8
12460 främjat 3
12461 främling 1
12462 främlingar 2
12463 främlingens 1
12464 främlings- 1
12465 främlingsfientlig 2
12466 främlingsfientliga 23
12467 främlingsfientlighet 25
12468 främlingsfientligheten 2
12469 främlingsfientlighetens 2
12470 främlingsfientligt 5
12471 främlingshat 1
12472 främlingsrädsla 1
12473 främlingsskap 1
12474 främmande 13
12475 främst 97
12476 främsta 39
12477 främste 2
12478 fräsanden 1
12479 fräsch 1
12480 fräste 1
12481 fråga 778
12482 frågade 24
12483 frågan 487
12484 frågande 6
12485 frågans 4
12486 frågar 50
12487 frågat 6
12488 frågekomplex 1
12489 frågeläge 5
12490 frågelägen 1
12491 frågelägesinställning 1
12492 frågeläget 1
12493 frågesatsen 1
12494 frågestunden 15
12495 frågeställaren 4
12496 frågeställningen 1
12497 frågetecken 4
12498 frågor 490
12499 frågorna 74
12500 från 1841
12501 frångår 1
12502 frånsett 1
12503 frånstötande 1
12504 frånsäga 1
12505 fråntar 1
12506 fråntas 3
12507 fråntog 1
12508 frånvarande 10
12509 frånvaro 8
12510 frånvaron 6
12511 frö 2
12512 fröet 1
12513 fröjdar 1
12514 fukt 1
12515 fuktigt 1
12516 full 69
12517 fulla 21
12518 fullare 1
12519 fullaste 1
12520 fullborda 2
12521 fullbordad 3
12522 fullbordandet 2
12523 fullbordar 1
12524 fullbordas 2
12525 fullbordat 1
12526 fullfölja 4
12527 fullföljas 1
12528 fullföljer 3
12529 fullföljt 1
12530 fullgjort 2
12531 fullgör 1
12532 fullgöra 7
12533 fullgöras 2
12534 fullgörs 1
12535 fullkomlig 1
12536 fullkomlighet 1
12537 fullkomligt 9
12538 fullkomnade 1
12539 fullmakt 2
12540 fullmaktsbestämmelser 1
12541 fullmäktige 1
12542 fullo 8
12543 fullpackad 1
12544 fullsatt 1
12545 fullständig 34
12546 fullständiga 10
12547 fullständigt 70
12548 fullt 62
12549 fulltecknade 1
12550 fulltoniga 1
12551 fullvärdig 6
12552 fullvärdiga 2
12553 fullända 1
12554 fulländar 1
12555 fulländat 1
12556 fult 1
12557 fumlig 1
12558 fundamental 1
12559 fundamentala 2
12560 fundamentalt 3
12561 fundera 18
12562 funderade 8
12563 funderar 8
12564 funderingar 3
12565 funderingarna 1
12566 fundersökningar 1
12567 fungera 56
12568 fungerade 2
12569 fungerande 23
12570 fungerar 58
12571 fungerat 8
12572 funktion 30
12573 funktionalistiska 2
12574 funktionella 1
12575 funktionellt 1
12576 funktionen 6
12577 funktioner 13
12578 funktionerna 4
12579 funktionsbrister 1
12580 funktionsduglig 1
12581 funktionsduglighet 3
12582 funktionshinder 8
12583 funktionsregler 2
12584 funktionssätt 1
12585 funktionsvillkor 1
12586 funktionärer 1
12587 funktionärers 1
12588 funnit 9
12589 funnits 23
12590 fusion 2
12591 fusionen 2
12592 fusioner 9
12593 fusionsförordningen 1
12594 fusionshaussen 1
12595 fusionskontrollen 1
12596 fusionsrätten 1
12597 fusk 1
12598 futtiga 2
12599 fylla 12
12600 fyllande 1
12601 fyllas 3
12602 fylld 2
12603 fyllda 2
12604 fyllde 5
12605 fylldes 1
12606 fyller 2
12607 fyllig 1
12608 fylls 1
12609 fyllt 7
12610 fyllts 2
12611 fyra 87
12612 fyrahundra 3
12613 fyratusen 1
12614 fyrkant 1
12615 fyrtio 8
12616 fyrtioett 1
12617 fyrtiosju 1
12618 fyrtiotalet 1
12619 fyrtioåtta 1
12620 fysiken 1
12621 fysiologiska 1
12622 fysisk 8
12623 fysiska 17
12624 fysiskt 7
12625 fädernearvet 1
12626 fällan 1
12627 fällde 2
12628 fäller 1
12629 fälls 1
12630 fällt 1
12631 fällts 3
12632 fält 37
12633 fältelement 1
12634 fälten 7
12635 fältet 19
12636 fältets 2
12637 fängelse 9
12638 fängelsedagbok 1
12639 fängelser 1
12640 fängelserna 3
12641 fängelsestraff 2
12642 fängslas 1
12643 fängslats 1
12644 färd 9
12645 färdades 1
12646 färdats 1
12647 färden 2
12648 färdig 4
12649 färdiga 2
12650 färdigheter 1
12651 färdigställa 1
12652 färdigställde 1
12653 färdigt 8
12654 färdriktning 1
12655 färg 3
12656 färgad 2
12657 färgade 2
12658 färgas 1
12659 färgen 4
12660 färger 6
12661 färgkombinationen 1
12662 färgskrubben 1
12663 färje- 1
12664 färjetrafiken 1
12665 färre 10
12666 färska 1
12667 färskt 2
12668 färskvatten 2
12669 färskvattenförsörjning 1
12670 fäst 3
12671 fästa 9
12672 fästad 1
12673 fästade 1
12674 fäste 1
12675 fäster 8
12676 fästning 1
12677 fästs 1
12678 få 650
12679 fåfänga 3
12680 fågel 3
12681 fågeldirektiven 1
12682 fågeldirektivet 1
12683 fågellivet 1
12684 fågelpopulationer 1
12685 fågelskrämma 1
12686 fågelskyddssällskapet 1
12687 fågelvänner 1
12688 fåglar 12
12689 fålla 1
12690 fån 1
12691 fånga 1
12692 fångade 3
12693 fångades 1
12694 fångar 13
12695 fångarna 6
12696 fångarnas 1
12697 fångars 1
12698 fångas 1
12699 fångat 3
12700 fånge 1
12701 fångna 2
12702 fångst 5
12703 fångsten 1
12704 fångster 2
12705 fångsterna 2
12706 fångstförbud 1
12707 fångstkvoter 1
12708 fångstmetoder 1
12709 fångstmängd 2
12710 fångstmängden 3
12711 får 575
12712 fårad 1
12713 fåret 1
12714 fårköttsproduktion 1
12715 fåror 1
12716 fås 2
12717 fåtal 10
12718 fåtalet 1
12719 fåtaliga 1
12720 fått 195
12721 fåtölj 1
12722 fåtöljer 1
12723 fåtöljerna 1
12724 föda 2
12725 födande 3
12726 född 2
12727 födda 3
12728 födde 1
12729 föddes 10
12730 födelse 1
12731 födelseakt 1
12732 födelsebygd 1
12733 födelsedag 1
12734 födelsedagen 1
12735 födelsedagskalasen 1
12736 födelseort 1
12737 födelsetal 1
12738 föder 4
12739 födoämnen 1
12740 föds 4
12741 födsel 2
12742 födseln 1
12743 föga 5
12744 följa 77
12745 följaktligen 36
12746 följande 111
12747 följas 12
12748 följd 67
12749 följde 17
12750 följden 5
12751 följder 14
12752 följderna 12
12753 följdes 5
12754 följdfråga 1
12755 följdfrågan 1
12756 följdfrågor 1
12757 följdriktig 1
12758 följdskador 1
12759 följdskadorna 1
12760 följdåtgärder 1
12761 följe 3
12762 följer 43
12763 följerätten 1
12764 följs 6
12765 följt 14
12766 följts 4
12767 föll 8
12768 fönster 7
12769 fönsterbrädan 1
12770 fönsterbrädet 1
12771 fönstergallret 1
12772 fönsterkarmar 1
12773 fönsterplats 1
12774 fönstren 3
12775 fönstret 14
12776 för 9583
12777 föra 81
12778 förakt 3
12779 föraktat 1
12780 föraktfull 1
12781 föraktfullt 1
12782 förankra 2
12783 förankrad 2
12784 förankrade 4
12785 förankras 1
12786 förankring 1
12787 föranleda 1
12788 föranledde 2
12789 föranleder 3
12790 föranslutningsavtal 1
12791 föranslutningsstrategi 2
12792 föranslutningsstrategin 3
12793 föranslutningsstöd 2
12794 förarbetet 1
12795 förare 2
12796 föraren 1
12797 förargat 1
12798 förargligt 1
12799 förarna 2
12800 föras 18
12801 förband 2
12802 förbannat 2
12803 förbannelse 2
12804 förbarmande 1
12805 förbaskat 1
12806 förbehåll 6
12807 förbehållas 3
12808 förbehållen 1
12809 förbehåller 2
12810 förbehållet 1
12811 förbehållslöst 1
12812 förbereda 20
12813 förberedande 14
12814 förberedandet 2
12815 förberedas 5
12816 förberedd 3
12817 förberedda 3
12818 förberedde 4
12819 förbereddes 1
12820 förberedelse 2
12821 förberedelse- 1
12822 förberedelsearbete 1
12823 förberedelsearbetet 1
12824 förberedelsen 2
12825 förberedelseperiod 1
12826 förberedelser 9
12827 förberedelserna 9
12828 förbereder 13
12829 förbereds 2
12830 förberett 4
12831 förberetts 2
12832 förbi 17
12833 förbifarten 2
12834 förbigå 1
12835 förbigående 9
12836 förbigår 1
12837 förbigås 2
12838 förbiilande 1
12839 förbinda 3
12840 förbindelse 14
12841 förbindelselänk 1
12842 förbindelsen 2
12843 förbindelser 39
12844 förbindelseramar 1
12845 förbindelserna 48
12846 förbindelsestrukturen 1
12847 förbinder 8
12848 förbindligheten 1
12849 förbiseende 2
12850 förbisprunget 1
12851 förbisprungits 1
12852 förbittrat 1
12853 förbittring 1
12854 förbjuda 13
12855 förbjudas 5
12856 förbjuden 2
12857 förbjuder 7
12858 förbjudet 7
12859 förbjudit 2
12860 förbjudna 4
12861 förbjuds 1
12862 förbjöd 1
12863 förbjöds 1
12864 förblev 1
12865 förbli 19
12866 förblir 23
12867 förblivande 1
12868 förblivit 1
12869 förbluffade 1
12870 förbluffande 1
12871 förbrukade 1
12872 förbrukar 1
12873 förbrukaren 1
12874 förbrukat 2
12875 förbrukning 2
12876 förbrukningen 1
12877 förbrukningsnivåer 1
12878 förbryllad 1
12879 förbryllande 1
12880 förbrytare 2
12881 förbrytelser 2
12882 förbrytelserna 1
12883 förbränning 1
12884 förbränningskvoten 1
12885 förbränns 1
12886 förbud 18
12887 förbudet 9
12888 förbudsförbehåll 1
12889 förbudsprincipen 1
12890 förbund 1
12891 förbunden 2
12892 förbundet 3
12893 förbundit 9
12894 förbundna 4
12895 förbundskansler 3
12896 förbundskanslern 1
12897 förbundsländer 1
12898 förbundsländerna 1
12899 förbundsregeringen 1
12900 förbundsrepubliken 1
12901 förbättra 105
12902 förbättrad 12
12903 förbättrade 6
12904 förbättrande 1
12905 förbättrar 12
12906 förbättras 19
12907 förbättrat 2
12908 förbättrats 9
12909 förbättring 31
12910 förbättringar 20
12911 förbättringen 4
12912 förbättringstendens 1
12913 förbättringsåtagande 1
12914 förda 3
12915 förde 15
12916 fördefinierade 2
12917 fördel 22
12918 fördela 3
12919 fördelad 1
12920 fördelade 3
12921 fördelaktigt 1
12922 fördelar 18
12923 fördelarna 7
12924 fördelas 7
12925 fördelat 3
12926 fördelats 1
12927 fördelen 4
12928 fördelning 15
12929 fördelningen 9
12930 fördelningsbegreppet 1
12931 fördelningsinstrument 1
12932 fördelningskriterierna 1
12933 fördelningsnyckel 1
12934 fördelningsnyckeln 1
12935 fördelningspolitik 2
12936 fördelningspolitiken 1
12937 fördes 3
12938 fördjupa 12
12939 fördjupad 4
12940 fördjupar 1
12941 fördjupas 2
12942 fördjupat 4
12943 fördjupning 4
12944 fördjupningen 2
12945 fördomar 2
12946 fördomsfrihet 1
12947 fördomsfullhet 1
12948 fördra 2
12949 fördrag 24
12950 fördragen 51
12951 fördragens 5
12952 fördraget 98
12953 fördragets 14
12954 fördrags 1
12955 fördragsanalfabeter 1
12956 fördragsartiklar 1
12957 fördragsfäst 1
12958 fördragsmässiga 1
12959 fördragsmässigt 1
12960 fördragsorganisationens 1
12961 fördragsreform 1
12962 fördragsreglerna 1
12963 fördragssituation 1
12964 fördragsslutande 2
12965 fördragstexten 1
12966 fördragstexterna 1
12967 fördragsändringar 2
12968 fördragsändringarna 1
12969 fördrev 1
12970 fördrivits 1
12971 fördrivna 1
12972 fördrivning 1
12973 fördröja 1
12974 fördröjas 1
12975 fördubbla 4
12976 fördubblade 1
12977 fördubblades 1
12978 fördubblas 1
12979 fördubbling 1
12980 fördunklat 1
12981 fördunklats 1
12982 fördämningar 1
12983 fördärva 3
12984 fördärvad 2
12985 fördärvat 1
12986 fördärvbringande 1
12987 fördärvlig 1
12988 fördöma 18
12989 fördömande 11
12990 fördömanden 2
12991 fördömandet 1
12992 fördömas 1
12993 fördömer 17
12994 fördömt 2
12995 fördömts 1
12996 före 100
12997 före-före 1
12998 förebild 9
12999 förebildsmodellen 1
13000 förebråelse 1
13001 förebråelser 1
13002 förebrående 1
13003 förebrås 2
13004 förebygga 18
13005 förebyggande 40
13006 förebyggandet 6
13007 förebyggas 2
13008 förebygger 1
13009 föredra 11
13010 föredrag 1
13011 föredragande 79
13012 föredraganden 158
13013 föredragandena 8
13014 föredragandenas 1
13015 föredragandens 25
13016 föredragandes 2
13017 föredragit 4
13018 föredragning 2
13019 föredragningslista 17
13020 föredragningslistan 101
13021 föredragningslistor 1
13022 föredragningslistorna 2
13023 föredrar 9
13024 föredrog 3
13025 föredöme 4
13026 föredömlig 1
13027 föredömliga 2
13028 föredömligt 4
13029 förefalla 1
13030 förefaller 45
13031 föreföll 4
13032 föregick 1
13033 föregiven 1
13034 föregripa 2
13035 föregripande 3
13036 föregriper 1
13037 föregripit 1
13038 föregå 2
13039 föregående 57
13040 föregångare 8
13041 föregångares 1
13042 föregångarna 1
13043 föregår 1
13044 föregås 1
13045 förehavanden 3
13046 förekom 3
13047 förekomma 14
13048 förekommande 10
13049 förekommas 1
13050 förekommer 32
13051 förekommit 12
13052 förekomsten 5
13053 förelegat 1
13054 föreligga 2
13055 föreliggande 17
13056 föreligger 29
13057 föreläsa 2
13058 föreläsning 1
13059 föreläsningen 1
13060 föreläste 1
13061 förelåg 1
13062 föremål 38
13063 föremålen 1
13064 föremålet 1
13065 fören 1
13066 förena 24
13067 förenad 2
13068 förenade 4
13069 förenar 4
13070 förenas 3
13071 förenat 1
13072 förenats 1
13073 förening 7
13074 föreningar 3
13075 föreningarna 1
13076 förenkla 9
13077 förenklad 1
13078 förenklade 4
13079 förenklande 1
13080 förenklar 3
13081 förenklas 1
13082 förenkling 6
13083 förenlig 4
13084 förenliga 7
13085 förenlighet 1
13086 förenligheten 1
13087 förenligt 4
13088 förenta 3
13089 föresats 1
13090 föresatsen 2
13091 föresatser 9
13092 föresatserna 1
13093 föresatt 1
13094 föresatte 1
13095 föreskrev 1
13096 föreskrift 2
13097 föreskrifter 16
13098 föreskrifterna 2
13099 föreskriva 6
13100 föreskrivande 2
13101 föreskriven 1
13102 föreskriver 19
13103 föreskrivit 1
13104 föreskrivits 3
13105 föreskrivna 1
13106 föreskrivs 12
13107 föreslagen 3
13108 föreslagit 40
13109 föreslagits 20
13110 föreslagna 43
13111 föreslog 16
13112 föreslogs 6
13113 föreslå 47
13114 föreslår 88
13115 föreslås 37
13116 förespegla 1
13117 förespeglar 1
13118 förespråka 6
13119 förespråkar 14
13120 förespråkare 6
13121 förespråkarna 2
13122 förespråkas 1
13123 förespråkat 2
13124 förespråkats 1
13125 föreställa 16
13126 föreställde 2
13127 föreställdes 1
13128 föreställer 5
13129 föreställning 1
13130 föreställningar 3
13131 föreställningar- 1
13132 föreställningen 1
13133 föreståeligt 1
13134 förestående 11
13135 föreståndare 1
13136 föresätter 1
13137 företa 3
13138 företag 211
13139 företagande 4
13140 företagaranda 9
13141 företagarandan 1
13142 företagare 12
13143 företagaren 2
13144 företagarna 7
13145 företagarorganisationer 1
13146 företagartillfällen 1
13147 företagarvärlden 1
13148 företagen 83
13149 företagens 32
13150 företaget 30
13151 företagets 4
13152 företags 3
13153 företags- 1
13154 företagsamhet 10
13155 företagsamma 1
13156 företagsandan 1
13157 företagsavtal 1
13158 företagsbeskattning 1
13159 företagsbeslutet 1
13160 företagsdemokratisering 1
13161 företagsekonomisk 1
13162 företagsekonomiska 3
13163 företagsekonomiskt 2
13164 företagsfusioner 1
13165 företagsförvärv 1
13166 företagsgrupper 2
13167 företagsgrupperna 2
13168 företagsinterna 1
13169 företagsjuristernas 2
13170 företagskoncentration 1
13171 företagskonsulter 1
13172 företagsledningen 1
13173 företagsledningens 2
13174 företagslikvidation 1
13175 företagslivet 1
13176 företagsnamn 1
13177 företagsnedläggning 1
13178 företagsnedläggningar 1
13179 företagspolitiken 1
13180 företagsråd 2
13181 företagsrådet 6
13182 företagsrådsdirektivet 1
13183 företagsskapande 1
13184 företagsstadgar 1
13185 företagsstruktur 1
13186 företagsstrukturen 2
13187 företagsstöd 2
13188 företagsstöden 1
13189 företagstalangen 1
13190 företagsutveckling 1
13191 företeelse 1
13192 företeelser 2
13193 företräda 7
13194 företrädandet 1
13195 företrädare 116
13196 företrädaren 4
13197 företrädares 3
13198 företrädarna 17
13199 företrädas 4
13200 företrädd 2
13201 företrädda 6
13202 företrädde 1
13203 företräde 5
13204 företräder 22
13205 företrädesvis 2
13206 företräds 3
13207 företrätt 1
13208 förevisas 1
13209 förevändning 7
13210 förevändningar 1
13211 förevändningen 2
13212 förfader 1
13213 förfall 2
13214 förfalla 1
13215 förfallit 1
13216 förfallna 2
13217 förfalskare 1
13218 förfalskas 5
13219 förfalskning 12
13220 förfalskningar 11
13221 förfalskningsutrustning 1
13222 förfarande 47
13223 förfarandefrågor 1
13224 förfaranden 32
13225 förfarandena 14
13226 förfarandet 46
13227 förfaringssätt 1
13228 förfasade 1
13229 förfasar 1
13230 författa 1
13231 författare 4
13232 författaren 3
13233 författares 1
13234 författarna 1
13235 författarnamnet 1
13236 författarnas 1
13237 författat 4
13238 författats 1
13239 författningar 1
13240 författningen 1
13241 författningsenliga 1
13242 författningsfrågor 1
13243 författningsrätt 1
13244 förfela 1
13245 förfiningsarbete 1
13246 förfjol 1
13247 förflutet 1
13248 förflutna 21
13249 förflutnas 1
13250 förflytta 5
13251 förflyttade 2
13252 förflyttar 2
13253 förflyttats 1
13254 förflyttning 6
13255 förflyttningar 1
13256 förflyttningen 1
13257 förfoga 8
13258 förfogande 31
13259 förfoganderätt 1
13260 förfogar 21
13261 förfront 2
13262 förfrysningsskador 1
13263 förfrågan 5
13264 förfrågningar 3
13265 förfäders 1
13266 förfäktar 1
13267 förfärande 5
13268 förfärlig 1
13269 förfärliga 3
13270 förfärligaste 1
13271 förfärligt 5
13272 förfång 3
13273 förfölja 2
13274 förföljare 1
13275 förföljda 1
13276 förföljde 2
13277 förföljelser 3
13278 förföljelserna 3
13279 förföljer 1
13280 förföljs 3
13281 förförisk 2
13282 förförnyelse 1
13283 förfört 1
13284 förgiftar 1
13285 förgiftning 2
13286 förgiftningen 1
13287 förglömma 2
13288 förglömmas 1
13289 förgrening 1
13290 förgrovande 1
13291 förgrunden 5
13292 förgät-mig-ej-blått 1
13293 förgäves 2
13294 förgångna 2
13295 förgångnas 1
13296 förhalande 1
13297 förhand 8
13298 förhandla 26
13299 förhandlade 1
13300 förhandlande 1
13301 förhandlar 3
13302 förhandlarna 2
13303 förhandlas 3
13304 förhandlat 2
13305 förhandlats 2
13306 förhandling 14
13307 förhandlingar 38
13308 förhandlingarna 54
13309 förhandlingarnas 1
13310 förhandlingen 15
13311 förhandlings- 2
13312 förhandlingsbordet 1
13313 förhandlingsflexibilitet 1
13314 förhandlingsforum 1
13315 förhandlingsförfarande 1
13316 förhandlingsgruppen 1
13317 förhandlingsklimatet 1
13318 förhandlingsmandatet 1
13319 förhandlingsparterna 1
13320 förhandlingspartnerna 1
13321 förhandlingsperiod 1
13322 förhandlingsposition 1
13323 förhandlingsprocess 2
13324 förhandlingsprocessen 3
13325 förhandlingsrunda 1
13326 förhandlingsrundan 3
13327 förhandlingsrundorna 1
13328 förhandlingssammanträde 1
13329 förhandlingssammanträdena 1
13330 förhandlingssammanträdet 1
13331 förhandlingssituation 1
13332 förhandlingsskicklighet 1
13333 förhandlingsärenden 1
13334 förhands- 1
13335 förhandsanmälningar 1
13336 förhandsavgörande 2
13337 förhandsavgöranden 1
13338 förhandsbekräftelse 1
13339 förhandsinformation 1
13340 förhandskontroll 2
13341 förhandskontrollen 2
13342 förhastade 3
13343 förhastar 1
13344 förhastat 2
13345 förhindra 72
13346 förhindrade 1
13347 förhindrande 1
13348 förhindrandet 1
13349 förhindrar 9
13350 förhindras 9
13351 förhindrat 2
13352 förhindrats 1
13353 förhistorisk 1
13354 förhoppning 8
13355 förhoppningar 18
13356 förhoppningen 7
13357 förhoppningsvis 8
13358 förhärskande 2
13359 förhålla 1
13360 förhållande 54
13361 förhållanden 45
13362 förhållandena 14
13363 förhållandet 30
13364 förhållandevis 3
13365 förhåller 7
13366 förhållit 1
13367 förhållningssätt 4
13368 förhållningssättet 2
13369 förhånas 1
13370 förhöjt 1
13371 förhöll 1
13372 förintas 1
13373 förintelse 1
13374 förintelsekonferensen 1
13375 förintelsen 1
13376 förirra 1
13377 förkasta 5
13378 förkastade 6
13379 förkastades 3
13380 förkastandet 1
13381 förkastar 8
13382 förkastas 2
13383 förkastat 1
13384 förkastats 2
13385 förkastligt 2
13386 förklara 34
13387 förklarade 23
13388 förklarar 93
13389 förklaras 9
13390 förklarat 11
13391 förklarats 5
13392 förklaring 19
13393 förklaringar 6
13394 förklaringarna 5
13395 förklaringen 4
13396 förklarliga 1
13397 förkläde 1
13398 förkläden 1
13399 förklädet 1
13400 förklädnad 1
13401 förknippad 2
13402 förknippade 5
13403 förknippas 1
13404 förkorta 3
13405 förkortad 1
13406 förkortade 3
13407 förkortas 2
13408 förkortat 1
13409 förkortning 1
13410 förkortningen 1
13411 förkovran 1
13412 förkromade 1
13413 förkrossande 1
13414 förkunna 1
13415 förkunnade 1
13416 förkunnar 1
13417 förkunnat 1
13418 förkunnats 1
13419 förkämpe 3
13420 förkänsla 1
13421 förlagen 1
13422 förlagor 2
13423 förledas 1
13424 förlegad 1
13425 förlegade 1
13426 förlika 1
13427 förlikar 1
13428 förlikning 13
13429 förlikningar 1
13430 förlikningen 13
13431 förliknings- 1
13432 förlikningsetappen 1
13433 förlikningsförfarande 5
13434 förlikningsförfarandet 9
13435 förlikningskommitté 1
13436 förlikningskommittén 11
13437 förlikningskommitténs 6
13438 förlikningsprocess 3
13439 förlikningsprocessen 2
13440 förlikningsvävnad 1
13441 förlisning 7
13442 förlisningen 3
13443 förliste 2
13444 förlita 8
13445 förlitar 8
13446 förloppet 1
13447 förlora 18
13448 förlorad 4
13449 förlorade 12
13450 förlorades 1
13451 förlorar 15
13452 förlorare 1
13453 förloras 1
13454 förlorat 28
13455 förlorats 1
13456 förlossningskliniker 1
13457 förlust 7
13458 förlustbringande 1
13459 förlusten 6
13460 förluster 13
13461 förlusterna 3
13462 förlutet 1
13463 förlägenhet 1
13464 förläggas 1
13465 förläggning 2
13466 förlänga 7
13467 förlängas 2
13468 förlängde 1
13469 förlänger 2
13470 förlängning 8
13471 förlängningen 4
13472 förlängs 4
13473 förlängts 2
13474 förlåt 1
13475 förlåta 2
13476 förlåten 1
13477 förlåter 1
13478 förlöjligar 1
13479 förlöper 1
13480 förmanad 1
13481 förmaning 1
13482 förmedla 9
13483 förmedlade 1
13484 förmedlande 1
13485 förmedlar 2
13486 förmedlare 1
13487 förmedlas 1
13488 förmedling 1
13489 förmenande 3
13490 förment 1
13491 förmenta 2
13492 förmiddag 8
13493 förmiddagen 3
13494 förmiddagens 2
13495 förmiddags 9
13496 förmildrande 1
13497 förmodade 1
13498 förmodar 7
13499 förmodas 1
13500 förmodligen 37
13501 förmyndarskap 1
13502 förmå 9
13503 förmåga 42
13504 förmågan 5
13505 förmån 44
13506 förmånen 1
13507 förmåner 6
13508 förmånligt 1
13509 förmånsavtalen 1
13510 förmånsbehandling 2
13511 förmånspaketet 1
13512 förmånstagare 1
13513 förmånstagarna 1
13514 förmånstillträde 1
13515 förmånsursprung 1
13516 förmår 2
13517 förmås 1
13518 förmått 3
13519 förmögen 1
13520 förmögna 1
13521 förmörkelsen 1
13522 förnamn 1
13523 förnedrande 2
13524 förnedring 1
13525 förneka 10
13526 förnekande 1
13527 förnekar 3
13528 förnekas 4
13529 förnekat 1
13530 förnuft 4
13531 förnuftet 4
13532 förnuftig 10
13533 förnuftiga 10
13534 förnuftigare 2
13535 förnuftigt 16
13536 förnufts- 1
13537 förnumstigt 1
13538 förnya 11
13539 förnyad 1
13540 förnyade 5
13541 förnyande 1
13542 förnyandet 1
13543 förnyar 1
13544 förnyas 2
13545 förnyat 1
13546 förnybar 8
13547 förnybara 40
13548 förnyelse 16
13549 förnyelsen 6
13550 förnyelseområden 1
13551 förnämlig 1
13552 förnämsta 2
13553 förnärma 1
13554 förnärmade 1
13555 förolämpande 2
13556 förolämpar 2
13557 förolämpas 1
13558 förolämpat 1
13559 förolämpning 3
13560 förorda 1
13561 förordar 5
13562 förordas 1
13563 förordna 1
13564 förordnanden 1
13565 förordnas 1
13566 förordning 85
13567 förordningar 15
13568 förordningarna 3
13569 förordningen 46
13570 förordningens 6
13571 förorena 2
13572 förorenad 1
13573 förorenade 3
13574 förorenande 10
13575 förorenar 19
13576 förorenare 2
13577 förorenaren 22
13578 förorenarens 3
13579 förorenarna 1
13580 förorenarnas 1
13581 förorenas 5
13582 förorenat 4
13583 förorenats 1
13584 förorening 15
13585 föroreningar 26
13586 föroreningarna 6
13587 föroreningarnas 1
13588 föroreningen 6
13589 föroreningsminskningar 1
13590 förorsaka 3
13591 förorsakad 1
13592 förorsakade 2
13593 förorsakar 2
13594 förorsakas 1
13595 förorsakat 3
13596 förorsakats 3
13597 förorter 5
13598 förorters 1
13599 förpackat 1
13600 förpackning 3
13601 förpackningar 1
13602 förpackningsdirektivet 1
13603 förpassa 2
13604 förpassade 1
13605 förpassades 1
13606 förpassas 1
13607 förpestade 1
13608 förpliktad 1
13609 förpliktade 3
13610 förpliktande 1
13611 förpliktar 3
13612 förpliktas 1
13613 förpliktelse 6
13614 förpliktelsen 3
13615 förpliktelser 14
13616 förpliktiga 1
13617 förpliktigad 2
13618 förpliktigade 2
13619 förpliktigande 1
13620 förpliktigar 1
13621 förpliktigas 1
13622 förpliktigat 3
13623 förr 15
13624 förra 118
13625 förre 6
13626 förresten 5
13627 förrgår 5
13628 förringa 2
13629 förringar 1
13630 förräderi 2
13631 förrädisk 1
13632 förrän 22
13633 förrättar 1
13634 förrättas 1
13635 förråd 1
13636 förrådde 1
13637 förs 18
13638 församlade 1
13639 församling 25
13640 församlingar 3
13641 församlingarna 2
13642 församlingen 27
13643 församlingens 2
13644 församlings 1
13645 försatt 2
13646 förse 18
13647 förseglad 1
13648 försena 4
13649 försenad 8
13650 försenade 7
13651 försenades 1
13652 försenar 1
13653 försenas 2
13654 försenat 5
13655 försening 7
13656 förseningar 8
13657 förseningarna 1
13658 förseningen 6
13659 förser 3
13660 förses 5
13661 försett 2
13662 försetts 1
13663 försiggick 1
13664 försiktig 7
13665 försiktiga 17
13666 försiktighet 14
13667 försiktigheten 2
13668 försiktighetsprincipen 58
13669 försiktighetsprinipen 1
13670 försiktighetsåtgärd 2
13671 försiktighetsåtgärden 1
13672 försiktighetsåtgärder 3
13673 försiktigt 7
13674 försjunken 1
13675 försjunket 1
13676 försjönk 1
13677 förskansad 1
13678 förskingra 1
13679 förskingrat 1
13680 förskingring 2
13681 förskjutas 1
13682 förskjutning 3
13683 förskolor 1
13684 förskonade 1
13685 förskottsbetalningar 1
13686 förskräcka 1
13687 förskräckande 1
13688 förskräcklig 2
13689 förskräckliga 1
13690 förskräckligt 1
13691 förskräckt 2
13692 förskräckta 1
13693 förslag 576
13694 förslagen 42
13695 förslaget 185
13696 förslagets 2
13697 förslagits 2
13698 förslagna 2
13699 förslagsdel 1
13700 förslagspaket 1
13701 förslagsstadiet 1
13702 förslagsställandet 1
13703 förslagsställaren 1
13704 förslavade 1
13705 förslår 2
13706 förslås 2
13707 förslösat 1
13708 försona 3
13709 försonande 3
13710 försoning 8
13711 försoningen 2
13712 försoningskommission 1
13713 försoningsprocessen 1
13714 försoningsprogrammet 2
13715 försonlig 1
13716 förspilla 1
13717 försprång 1
13718 först 140
13719 första 579
13720 förstabehandling 1
13721 förstabehandlingen 2
13722 förstainstansrätt 2
13723 förstainstansrätten 16
13724 förstainstansrättens 3
13725 förstaklasspelare 1
13726 förste 3
13727 förstesekreteraren 1
13728 förstfödde 1
13729 förstklassigt 1
13730 förstnämndas 1
13731 förstod 15
13732 förströdd 1
13733 förstulet 1
13734 förställer 1
13735 förställningskonsten 1
13736 förstärka 31
13737 förstärkande 1
13738 förstärkas 7
13739 förstärker 2
13740 förstärkning 15
13741 förstärks 7
13742 förstärkt 11
13743 förstärkta 3
13744 förstå 58
13745 förståeliga 1
13746 förståeligt 5
13747 förståelse 27
13748 förståelsen 2
13749 förstånd 1
13750 förståndiga 2
13751 förstår 71
13752 förstås 21
13753 förstått 22
13754 förstör 18
13755 förstöra 7
13756 förstöras 3
13757 förstörd 1
13758 förstörda 3
13759 förstörde 1
13760 förstördes 4
13761 förstörelse 5
13762 förstörelsen 7
13763 förstöringen 1
13764 förstörs 7
13765 förstört 3
13766 förstörts 8
13767 försumbar 1
13768 försumlighet 1
13769 försumma 1
13770 försummade 1
13771 försummar 2
13772 försummas 1
13773 försummat 1
13774 försummelse 4
13775 försummelsen 1
13776 försummelser 2
13777 försvaga 8
13778 försvagad 1
13779 försvagade 3
13780 försvagades 1
13781 försvagar 7
13782 försvagas 7
13783 försvagats 2
13784 försvagning 3
13785 försvann 11
13786 försvar 31
13787 försvara 43
13788 försvarade 4
13789 försvarades 1
13790 försvarar 18
13791 försvarare 6
13792 försvaras 6
13793 försvarat 10
13794 försvarbara 2
13795 försvaret 11
13796 försvarets 1
13797 försvars- 2
13798 försvarsadvokat 1
13799 försvarsanslag 1
13800 försvarsbeslut 1
13801 försvarsbesparingar 1
13802 försvarsbudgetarna 1
13803 försvarsbudgeten 1
13804 försvarsfrågor 2
13805 försvarshållningen 1
13806 försvarsidentitet 2
13807 försvarsidentiteten 2
13808 försvarsindustrin 1
13809 försvarsinstinkt 1
13810 försvarskapacitet 1
13811 försvarskapaciteten 1
13812 försvarskostnader 1
13813 försvarslösa 2
13814 försvarsmaktens 1
13815 försvarsmedel 1
13816 försvarsminister 2
13817 försvarsministermöte 1
13818 försvarsministern 3
13819 försvarsministrarna 2
13820 försvarsministrarnas 1
13821 försvarsområdet 1
13822 försvarspolitik 18
13823 försvarspolitiken 6
13824 försvarsstrukturer 1
13825 försvarsstyrkor 1
13826 försvarsuppgifter 1
13827 försvarsuppgifterna 1
13828 försvarsutgifter 2
13829 försvarsutvecklingsarbete 1
13830 försvinna 10
13831 försvinnande 2
13832 försvinner 30
13833 försvunnen 1
13834 försvunnit 9
13835 försvåra 2
13836 försvårande 1
13837 försvårar 3
13838 försvåras 3
13839 försäkra 40
13840 försäkrade 6
13841 försäkran 2
13842 försäkrar 7
13843 försäkrats 1
13844 försäkring 1
13845 försäkringar 9
13846 försäkringarna 1
13847 försäkringsavgifter 1
13848 försäkringsbedrägerier 1
13849 försäkringsbevis 3
13850 försäkringsbolag 2
13851 försäkringsbolagen 1
13852 försäkringsbolaget 1
13853 försäkringsmarknaden 1
13854 försäkringsrättigheter 1
13855 försäkringssektorn 1
13856 försäkringsskydd 2
13857 försäkringssystem 1
13858 försäkringssystemen 1
13859 försäljaren 2
13860 försäljning 8
13861 försäljningen 2
13862 försäljningsnedgången 2
13863 försäljningsrapport 1
13864 försäljningsrapporten 1
13865 försäljningsvolym 1
13866 försäljs 1
13867 försämra 5
13868 försämrad 3
13869 försämrade 4
13870 försämrande 1
13871 försämras 6
13872 försämring 4
13873 försämringar 1
13874 försämringarna 1
13875 försämringen 3
13876 försändelserna 1
13877 försänkts 1
13878 försätter 1
13879 försåg 2
13880 försågs 1
13881 försåtligt 1
13882 försåvitt 1
13883 försök 30
13884 försöka 108
13885 försöken 4
13886 försöker 75
13887 försöket 3
13888 försökslaboratorium 1
13889 försöksmässigt 1
13890 försökt 23
13891 försökte 37
13892 försökts 1
13893 försörja 3
13894 försörjer 1
13895 försörjning 4
13896 försörjningsgrund 1
13897 fört 13
13898 förtal 1
13899 förtecken 1
13900 förtecknades 1
13901 förteckning 7
13902 förteckningen 7
13903 förtid 1
13904 förtida 1
13905 förtidspension 2
13906 förtidspensionerade 2
13907 förtidspensionering 2
13908 förtidspensioneringssystemet 2
13909 förtjusande 1
13910 förtjusning 3
13911 förtjust 4
13912 förtjusta 2
13913 förtjäna 4
13914 förtjänade 2
13915 förtjänar 40
13916 förtjänats 1
13917 förtjänst 2
13918 förtjänsten 2
13919 förtjänster 3
13920 förtjänstfulla 1
13921 förtjänstfullt 2
13922 förtjänt 1
13923 förtjänta 2
13924 förtroende 67
13925 förtroendeförskott 1
13926 förtroendeklyftan 1
13927 förtroendekris 2
13928 förtroendeposter 1
13929 förtroenderöst 1
13930 förtroendeskapande 3
13931 förtroendet 17
13932 förtroendeuppbyggnaden 1
13933 förtroendevald 4
13934 förtroendevalda 2
13935 förtroendeväckande 1
13936 förtrogen 1
13937 förtrogna 1
13938 förtrollar 1
13939 förtrollat 1
13940 förtryck 4
13941 förtryckande 2
13942 förtryckare 1
13943 förtryckarhierarki 1
13944 förtryckarregimen 1
13945 förtrycket 2
13946 förtrycktas 1
13947 förtrytelse 1
13948 förträffliga 2
13949 förträfflighet 1
13950 förtränger 1
13951 förts 11
13952 förtursbehandling 1
13953 förtvivla 1
13954 förtvivlade 3
13955 förtvivlan 5
13956 förtvivlat 2
13957 förtydliga 6
13958 förtydligande 2
13959 förtydliganden 4
13960 förtäckt 2
13961 förtäckta 2
13962 förtära 1
13963 förtärande 1
13964 förtätad 1
13965 förtöjd 1
13966 förtöjda 1
13967 förunderligt 2
13968 förundersökningshandlingar 1
13969 förundra 1
13970 förut 11
13971 förutan 1
13972 förutbestämd 1
13973 förutbestämt 1
13974 förutom 42
13975 förutsatt 3
13976 förutsatte 1
13977 förutse 6
13978 förutsebar 1
13979 förutsedd 1
13980 förutseende 2
13981 förutser 1
13982 förutses 5
13983 förutsett 2
13984 förutsetts 3
13985 förutspå 1
13986 förutspåddes 2
13987 förutspås 1
13988 förutsäga 3
13989 förutsägbar 2
13990 förutsägbara 1
13991 förutsägbart 1
13992 förutsägelse 1
13993 förutsätta 2
13994 förutsättas 1
13995 förutsätter 30
13996 förutsättning 39
13997 förutsättningar 24
13998 förutsättningarna 11
13999 förutsättningen 4
14000 förutsättningslös 1
14001 förutsätts 1
14002 förutvarande 3
14003 förvalta 11
14004 förvaltad 2
14005 förvaltande 1
14006 förvaltar 4
14007 förvaltare 2
14008 förvaltaren 2
14009 förvaltas 4
14010 förvaltning 62
14011 förvaltningar 6
14012 förvaltningarna 2
14013 förvaltningarnas 1
14014 förvaltningen 36
14015 förvaltningens 1
14016 förvaltningsbolag 6
14017 förvaltningsbolagen 3
14018 förvaltningsbolaget 1
14019 förvaltningsförfarande 3
14020 förvaltningsförfaranden 1
14021 förvaltningsförfarandet 3
14022 förvaltningskommittéer 1
14023 förvaltningskostnaderna 2
14024 förvaltningsmyndigheters 1
14025 förvaltningsområde 1
14026 förvaltningsorgan 1
14027 förvaltningsprinciper 1
14028 förvaltningsrätt 2
14029 förvaltningssed 1
14030 förvaltningsstrukturen 1
14031 förvaltningssystem 3
14032 förvaltningstekniska 1
14033 förvaltningsuppdrag 1
14034 förvaltningsuppgifterna 1
14035 förvaltningsverksamhet 1
14036 förvaltningsåtgärder 1
14037 förvaltningsåtgärderna 1
14038 förvandla 6
14039 förvandlade 1
14040 förvandlar 5
14041 förvandlas 8
14042 förvandlat 1
14043 förvandlats 4
14044 förvanskar 1
14045 förvanskas 1
14046 förvanskats 1
14047 förvar 1
14048 förvaras 1
14049 förvarna 1
14050 förvarnade 1
14051 förvarningssystem 1
14052 förverkliga 23
14053 förverkligades 1
14054 förverkligande 1
14055 förverkligandet 6
14056 förverkligas 13
14057 förverkligats 4
14058 förvirrad 3
14059 förvirrade 1
14060 förvirrande 2
14061 förvirrar 1
14062 förvirrat 2
14063 förvirring 12
14064 förvirringen 1
14065 förvisade 1
14066 förvisats 1
14067 förvisningsorder 1
14068 förvissad 2
14069 förvissade 1
14070 förvissning 1
14071 förvisso 22
14072 förvriden 1
14073 förvränga 1
14074 förvrängd 1
14075 förväg 21
14076 förvägra 2
14077 förvägrad 1
14078 förvägrades 2
14079 förvägrar 2
14080 förvägras 1
14081 förvägrats 2
14082 förvänta 9
14083 förväntade 2
14084 förväntades 2
14085 förväntan 2
14086 förväntar 45
14087 förväntas 7
14088 förväntat 4
14089 förväntningar 18
14090 förväntningarna 5
14091 förvärra 2
14092 förvärrade 1
14093 förvärras 5
14094 förvärrat 2
14095 förvärrats 3
14096 förvärva 4
14097 förvärvas 1
14098 förvärvat 1
14099 förvärvsarbete 4
14100 förvärvsarbetet 2
14101 förväxla 2
14102 förväxlar 1
14103 förvåna 2
14104 förvånad 6
14105 förvånade 3
14106 förvånande 3
14107 förvånansvärt 3
14108 förvånar 2
14109 förvånas 2
14110 förvånats 1
14111 förvåning 3
14112 förädla 2
14113 förädlade 2
14114 förälder 1
14115 föräldraledighet 2
14116 föräldrar 15
14117 föräldrarnas 1
14118 föräldrars 3
14119 förälskad 1
14120 föränderliga 2
14121 förändra 27
14122 förändrade 4
14123 förändrades 3
14124 förändrar 5
14125 förändras 21
14126 förändrat 3
14127 förändrats 8
14128 förändring 42
14129 förändringar 65
14130 förändringarna 12
14131 förändringen 3
14132 förändringens 1
14133 förändringsarbetet 2
14134 förändringsprocesser 1
14135 föråldrad 1
14136 föråldrade 10
14137 föråldrat 2
14138 förödande 11
14139 förödelse 3
14140 förödmjukande 1
14141 förödmjukelser 1
14142 förökar 1
14143 förökning 1
14144 förövades 1
14145 förövaren 2
14146 förövarna 2
14147 föröver 1
14148 fötter 8
14149 fötterna 6
14150 fötts 2
14151 g 3
14152 gaffel 3
14153 gaffeldukar 1
14154 gaffeln 1
14155 gafflarnas 1
14156 gagn 4
14157 gagna 1
14158 gagnar 3
14159 gagnat 2
14160 galakvinnor 1
14161 galax 1
14162 galaxer 1
14163 galen 4
14164 galenskapen 1
14165 galenskaps 1
14166 galiciska 1
14167 galjonsfiguren 1
14168 galleon 1
14169 galler 1
14170 gallerstängerna 2
14171 gallret 2
14172 gallringen 1
14173 galna 5
14174 galningar 1
14175 galopp 1
14176 gamla 87
14177 gamle 3
14178 gammal 22
14179 gammaldags 1
14180 gammalmodig 1
14181 gammalt 7
14182 gangstertyper 1
14183 ganska 87
14184 gapade 1
14185 gapet 1
14186 gapskratt 2
14187 garage 1
14188 garant 6
14189 garantera 116
14190 garanterad 2
14191 garanterade 4
14192 garanterar 31
14193 garanteras 13
14194 garanterat 6
14195 garanterats 1
14196 garanti 19
14197 garantier 30
14198 garantierna 9
14199 garantifonden 3
14200 garantin 5
14201 garantisektion 1
14202 garantisektionen 1
14203 garantisystemet 1
14204 garde-länderna 2
14205 garderobsdörren 1
14206 gardinen 1
14207 garn 1
14208 gas 1
14209 gaskammare 1
14210 gassade 1
14211 gasutsläpp 1
14212 gata 2
14213 gatan 24
14214 gathörn 1
14215 gathörnstyper 1
14216 gator 4
14217 gatorna 6
14218 gatornas 1
14219 gav 68
14220 gavel 2
14221 gavs 10
14222 ge 403
14223 gedigen 1
14224 gediget 1
14225 gedigna 2
14226 gehör 2
14227 gelikar 1
14228 gemener 3
14229 gemensam 140
14230 gemensamma 388
14231 gemensamt 57
14232 gemenskap 23
14233 gemenskapen 129
14234 gemenskapens 184
14235 gemenskaper 1
14236 gemenskaperna 5
14237 gemenskapernas 8
14238 gemenskaplig 1
14239 gemenskaps- 1
14240 gemenskapsarvet 1
14241 gemenskapsaspekt 1
14242 gemenskapsavtal 1
14243 gemenskapsbefogenheterna 1
14244 gemenskapsbestämmelser 2
14245 gemenskapsbestämmelserna 3
14246 gemenskapsbidrag 1
14247 gemenskapsbidraget 1
14248 gemenskapsbudgeten 5
14249 gemenskapsdimensionen 1
14250 gemenskapsdirektiv 2
14251 gemenskapsdirektiven 2
14252 gemenskapsengagemang 1
14253 gemenskapsfilosofin 1
14254 gemenskapsfond 2
14255 gemenskapsfonder 1
14256 gemenskapsfrågor 1
14257 gemenskapsfördragens 1
14258 gemenskapsgrupper 2
14259 gemenskapshamnar 1
14260 gemenskapshamnarna 1
14261 gemenskapshamnarnas 1
14262 gemenskapsinförlivande 1
14263 gemenskapsinitiativ 20
14264 gemenskapsinitiativen 13
14265 gemenskapsinitiativet 26
14266 gemenskapsinitiativets 1
14267 gemenskapsinitiativs 1
14268 gemenskapsinsatserna 1
14269 gemenskapsinstitutionerna 4
14270 gemenskapsinstitutionernas 3
14271 gemenskapsinstrument 3
14272 gemenskapsintresse 1
14273 gemenskapsintressen 1
14274 gemenskapskonstruktion 1
14275 gemenskapskontroll 1
14276 gemenskapslag 1
14277 gemenskapslagstiftning 5
14278 gemenskapslagstiftningen 13
14279 gemenskapslagstiftningens 1
14280 gemenskapsmaskinen 1
14281 gemenskapsmaskinens 1
14282 gemenskapsmedborgare 1
14283 gemenskapsnivå 28
14284 gemenskapsnormerna 1
14285 gemenskapsområdet 1
14286 gemenskapsorgan 2
14287 gemenskapspelaren 3
14288 gemenskapsplanet 1
14289 gemenskapspolitik 5
14290 gemenskapspolitiken 6
14291 gemenskapspolitikens 2
14292 gemenskapspreferensen 1
14293 gemenskapsprocessen 1
14294 gemenskapsproduktionen 1
14295 gemenskapsprogram 5
14296 gemenskapsprogrammen 5
14297 gemenskapsprogrammet 1
14298 gemenskapsram 2
14299 gemenskapsramen 1
14300 gemenskapsregister 1
14301 gemenskapsregler 2
14302 gemenskapsreglerna 5
14303 gemenskapsresurserna 2
14304 gemenskapsrätt 1
14305 gemenskapsrätten 17
14306 gemenskapsstadga 1
14307 gemenskapsstrategi 1
14308 gemenskapsstrukturerna 1
14309 gemenskapsstöd 2
14310 gemenskapsstödets 1
14311 gemenskapsstödramar 1
14312 gemenskapsstödramarna 1
14313 gemenskapsstödramen 11
14314 gemenskapssystem 1
14315 gemenskapstexter 1
14316 gemenskapsvatten 2
14317 gemenskapsvattnen 1
14318 gemenskapsåtgärd 1
14319 gemenskapsåtgärder 6
14320 gement 1
14321 gemyt 1
14322 gemål 1
14323 genant 1
14324 genast 24
14325 gender 7
14326 genderkurser 1
14327 genderutbildning 1
14328 genderutbildningen 1
14329 genera 1
14330 generad 3
14331 generade 1
14332 general 4
14333 generaladvokaten 1
14334 generalangrepp 1
14335 generaldirektorat 10
14336 generaldirektoraten 3
14337 generaldirektoratet 9
14338 generaldirektör 2
14339 generaldirektören 1
14340 generaldirektörens 1
14341 generaler 1
14342 generalförsamling 1
14343 generalförsamlingen 2
14344 generalisera 1
14345 generaliserade 1
14346 generaliseras 1
14347 generaliseringar 1
14348 generalklausul 1
14349 generalsekretariat 1
14350 generalsekreterare 22
14351 generalsekreteraren 3
14352 generalsekreterares 2
14353 generande 2
14354 generation 2
14355 generationen 2
14356 generationer 11
14357 generationerna 2
14358 generationernas 2
14359 generationers 1
14360 generell 8
14361 generella 9
14362 generellt 12
14363 generera 3
14364 genererar 7
14365 genereras 1
14366 generiska 1
14367 generositet 3
14368 generositeten 1
14369 generös 4
14370 generösa 1
14371 generösare 1
14372 generöst 3
14373 genetiskt 25
14374 gengäld 4
14375 gengångare 1
14376 genial 1
14377 genljud 1
14378 genmodifieringsteknik 1
14379 genom 678
14380 genomarbetad 1
14381 genomarbetat 2
14382 genomblickbar 2
14383 genomblickbarhet 5
14384 genomblickbarheten 1
14385 genomblickbart 3
14386 genomblåstes 1
14387 genombrott 5
14388 genombrottet 1
14389 genomdriva 6
14390 genomdrivande 1
14391 genomdrivit 1
14392 genomdrivs 2
14393 genomfarter 1
14394 genomför 18
14395 genomföra 144
14396 genomförande 34
14397 genomförandebefogenheter 4
14398 genomförandebeslut 1
14399 genomförandebestämmelserna 1
14400 genomföranden 1
14401 genomförandena 1
14402 genomförandet 76
14403 genomförandeverksamheterna 1
14404 genomförandeåtgärd 1
14405 genomförandeåtgärden 2
14406 genomförandeåtgärder 3
14407 genomföras 55
14408 genomförbar 5
14409 genomförbara 4
14410 genomförbarhet 2
14411 genomförbarheten 1
14412 genomförbart 4
14413 genomförd 4
14414 genomförda 3
14415 genomförde 5
14416 genomfördes 9
14417 genomförs 39
14418 genomfört 8
14419 genomförts 18
14420 genomgick 3
14421 genomgripande 16
14422 genomgå 5
14423 genomgående 3
14424 genomgång 4
14425 genomgången 1
14426 genomgår 5
14427 genomgått 7
14428 genomled 1
14429 genomlidandet 1
14430 genomläsning 3
14431 genomskinliga 2
14432 genomskinligt 1
14433 genomslag 4
14434 genomslagskraft 2
14435 genomsnitt 12
14436 genomsnittet 6
14437 genomsnittlig 4
14438 genomsnittliga 5
14439 genomsnittligen 1
14440 genomsnittligt 1
14441 genomsnittsregionerna 1
14442 genomströmmar 1
14443 genomsynlighet 1
14444 genomsyra 4
14445 genomsyrade 1
14446 genomsyrar 1
14447 genomsyras 2
14448 genomsyrats 1
14449 genomsöks 1
14450 genomsökte 1
14451 genomträngande 2
14452 genomträngning 1
14453 genomtänkt 1
14454 genomtänkta 1
14455 gensvar 2
14456 gentemot 78
14457 gentjänster 1
14458 genuin 2
14459 genusdimensionen 1
14460 geografisk 5
14461 geografiska 20
14462 geografiskt 5
14463 geologiska 1
14464 geologiskt 1
14465 geometri 1
14466 geopolitiska 2
14467 geostrategiska 3
14468 geostrategiskt 1
14469 ger 217
14470 ges 46
14471 gest 11
14472 gestalt 1
14473 gestalta 1
14474 gester 1
14475 gesterna 1
14476 gestikulerade 1
14477 gestikulerande 1
14478 geting 1
14479 gett 67
14480 getter 2
14481 getton 2
14482 getts 2
14483 gevär 1
14484 geväret 1
14485 ghananer 1
14486 ghetto 1
14487 gick 108
14488 gift 2
14489 gifta 2
14490 giftblandningarna 1
14491 gifte 3
14492 giftig 1
14493 giftiga 6
14494 giftigt 1
14495 giftkatastrof 1
14496 giftutsläppet 1
14497 gigantisk 2
14498 gigantiska 4
14499 gigantiskt 1
14500 giljotinen 1
14501 gilla 3
14502 gillade 1
14503 gillades 1
14504 gillande 3
14505 gillar 4
14506 gillrat 1
14507 giltig 5
14508 giltiga 2
14509 giltighet 6
14510 giltigheten 3
14511 giltighetstid 11
14512 giltighetstiden 3
14513 giltigt 3
14514 gin 2
14515 ginge 1
14516 giromedel 1
14517 gissa 4
14518 gissade 1
14519 gisslan 4
14520 gitarrer 1
14521 givande 3
14522 givandet 1
14523 givare 9
14524 givares 1
14525 givarkonferensen 1
14526 givarlandens 1
14527 givarlandet 1
14528 givarländer 1
14529 givarländerna 2
14530 givarna 6
14531 givarnas 1
14532 givarsamfundet 1
14533 givas 1
14534 given 2
14535 gives 1
14536 givet 3
14537 givetvis 72
14538 givit 12
14539 givits 2
14540 givmild 1
14541 givna 3
14542 gjord 2
14543 gjorda 1
14544 gjorde 108
14545 gjordes 16
14546 gjort 203
14547 gjorts 56
14548 glad 54
14549 glada 7
14550 gladde 2
14551 gladeligen 1
14552 glans 2
14553 glansdager 1
14554 glas 9
14555 glasdörr 1
14556 glasen 1
14557 glaset 1
14558 glashus 1
14559 glasklart 1
14560 glasmonter 1
14561 glasmontrarna 1
14562 glaspärlor 1
14563 glass 1
14564 glassförsäljarnas 1
14565 glasskivorna 1
14566 glasögon 3
14567 glasögonbärare 1
14568 glasögonen 3
14569 glatt 4
14570 gled 5
14571 glesa 1
14572 glesbefolkade 3
14573 glesbygden 1
14574 glesbygdsområden 1
14575 glest 3
14576 glida 1
14577 glider 2
14578 glimma 1
14579 glimmade 3
14580 glimmande 1
14581 glimmar 1
14582 glimt 1
14583 glimtar 1
14584 glitterögd 1
14585 glittrande 2
14586 global 17
14587 globala 30
14588 globaliserad 3
14589 globaliserade 4
14590 globaliserande 1
14591 globalisering 12
14592 globaliseringen 32
14593 globaliseringens 3
14594 globaliseringsdiskussionen 1
14595 globaliseringsprocessen 1
14596 globaliteten 1
14597 globalt 13
14598 glodde 1
14599 glorifiering 1
14600 glunkades 1
14601 glupskhet 1
14602 gläder 58
14603 glädja 14
14604 glädjande 15
14605 glädjas 4
14606 glädje 17
14607 glädjen 1
14608 glädjevitt 1
14609 gläds 12
14610 glänsande 3
14611 glänste 1
14612 glöd 2
14613 glödhög 1
14614 glödlampa 1
14615 glödlampor 1
14616 glöm 1
14617 glömde 6
14618 glömma 44
14619 glömmas 1
14620 glömmer 10
14621 glöms 1
14622 glömska 1
14623 glömskan 1
14624 glömt 9
14625 gnista 1
14626 gnistor 1
14627 gnistrade 1
14628 gnistrande 1
14629 gnistregnet 1
14630 gnuggar 1
14631 gnutta 2
14632 gnället 1
14633 goals 2
14634 god 65
14635 goda 94
14636 godafton 1
14637 godas 1
14638 gode 1
14639 godhjärtad 1
14640 godkänd 5
14641 godkända 8
14642 godkände 19
14643 godkändes 11
14644 godkänna 49
14645 godkännande 30
14646 godkännandeförbehåll 1
14647 godkännandena 1
14648 godkännandet 9
14649 godkännas 18
14650 godkänner 29
14651 godkänns 4
14652 godkänt 21
14653 godkänts 22
14654 godmodigt 1
14655 godo 5
14656 gods 39
14657 godset 1
14658 godsets 1
14659 godsfinka 1
14660 godstransporter 1
14661 godstransporterna 1
14662 godta 23
14663 godtagbar 9
14664 godtagbara 7
14665 godtagbart 17
14666 godtagit 3
14667 godtagits 1
14668 godtar 15
14669 godtas 11
14670 godtog 4
14671 godtogs 3
14672 godtycke 1
14673 godtycklig 2
14674 godtyckliga 2
14675 godtyckligt 4
14676 gojernas 1
14677 golfförsäljningen 2
14678 golvet 3
14679 gom 1
14680 good 3
14681 gossarna 1
14682 gosse 1
14683 gossen 1
14684 gott 48
14685 gottgöra 2
14686 gottgörelse 1
14687 gottgörelsen 1
14688 governance 5
14689 government 1
14690 governments 1
14691 governo 2
14692 grabb 1
14693 gracila 1
14694 graciös 1
14695 grad 61
14696 graden 5
14697 grader 9
14698 graderna 1
14699 gradvis 16
14700 gradvisa 4
14701 gradvist 1
14702 graecas 1
14703 grafiskt 1
14704 gram 4
14705 grammofonnål 1
14706 grammofonskivor 1
14707 granadillpuddingen 1
14708 granaterna 1
14709 grand 6
14710 grannar 12
14711 granne 1
14712 grannförbindelser 1
14713 grannlagenhet 1
14714 grannland 1
14715 grannlandet 2
14716 grannländer 4
14717 grannländerna 9
14718 grannländernas 1
14719 grannregioner 1
14720 grannregionernas 1
14721 grannskap 2
14722 grannskapet 2
14723 grannsämja 1
14724 grannsämjan 1
14725 granska 44
14726 granskade 7
14727 granskades 1
14728 granskar 8
14729 granskas 14
14730 granskat 3
14731 granskats 3
14732 granskning 31
14733 granskningar 1
14734 granskningarna 2
14735 granskningen 9
14736 granskningsenhet 1
14737 granskningsmekanismer 1
14738 granskningsprocess 3
14739 granskningssystemet 1
14740 gras 1
14741 gras-fest 1
14742 gras-fester 1
14743 gratis 12
14744 gratulationer 8
14745 gratulera 64
14746 gratulerade 1
14747 gratulerar 21
14748 gratulerat 1
14749 grav 3
14750 grava 1
14751 gravar 3
14752 graverande 4
14753 gravgrottor 1
14754 gravida 3
14755 graviditet 1
14756 gravt 1
14757 gravvalv 1
14758 green 1
14759 grejor 1
14760 grek 1
14761 grekcypriotiska 2
14762 grekerna 2
14763 grekisk-turkiska 1
14764 grekiska 28
14765 grekiskt 1
14766 gren 2
14767 grenar 3
14768 grenarna 2
14769 grenen 2
14770 grep 2
14771 grepen 1
14772 grepp 5
14773 greppa 1
14774 greppade 1
14775 greps 2
14776 grevskapsrådet 1
14777 grillad 1
14778 grillade 1
14779 grimas 2
14780 grimaserande 1
14781 grimskaft 2
14782 grina 1
14783 gripa 6
14784 gripas 1
14785 griper 3
14786 gripit 2
14787 gripna 1
14788 grips 1
14789 grisfet 1
14790 grissinistänger 1
14791 grogrund 1
14792 grogrunden 1
14793 grop 2
14794 groteska 1
14795 group 1
14796 grov 1
14797 grova 1
14798 grund 316
14799 grund- 2
14800 grunda 2
14801 grundad 11
14802 grundade 4
14803 grundades 4
14804 grundandet 2
14805 grundar 24
14806 grundarna 2
14807 grundas 13
14808 grundat 14
14809 grundbegrepp 1
14810 grundbulten 1
14811 grunddokument 2
14812 grunden 60
14813 grundens 1
14814 grunder 13
14815 grunderna 3
14816 grundfördrag 1
14817 grundförståelsen 1
14818 grundförtroende 1
14819 grundförutsättning 2
14820 grundförutsättningar 1
14821 grundidén 1
14822 grundingredienserna 1
14823 grundinställning 2
14824 grundkoncept 2
14825 grundkurs 1
14826 grundlagsstridigt 1
14827 grundlig 6
14828 grundliga 4
14829 grundligare 2
14830 grundligt 13
14831 grundläggande 238
14832 grundläggarna 1
14833 grundorsakerna 1
14834 grundpelare 1
14835 grundpelaren 1
14836 grundprincip 2
14837 grundprincipen 2
14838 grundprinciper 1
14839 grundprinciperna 2
14840 grundproblem 1
14841 grundproblemet 1
14842 grundregeln 1
14843 grundsatsen 3
14844 grundsatserna 1
14845 grundskolan 1
14846 grundskolebarn 1
14847 grundskolorna 1
14848 grundsten 2
14849 grundstenar 1
14850 grundstomme 1
14851 grundstommen 2
14852 grundsyn 1
14853 grundtankarna 1
14854 grundtes 1
14855 grundtonen 1
14856 grundtrygghet 1
14857 grundtryggheten 1
14858 grundutbildning 2
14859 grundval 52
14860 grundvalar 3
14861 grundvalen 2
14862 grundvatten 5
14863 grundvattenakviferer 1
14864 grundvattenförekomsternas 1
14865 grundvattenkvalitet 1
14866 grundvattenkvaliteten 1
14867 grundvattenlagren 1
14868 grundvattenreserverna 2
14869 grundvattenstatus 2
14870 grundvattenstatusen 1
14871 grundvattnet 11
14872 grundvillkor 1
14873 grundämnen 1
14874 grupp 221
14875 gruppen 67
14876 gruppens 10
14877 grupper 78
14878 gruppera 2
14879 grupperade 3
14880 grupperas 1
14881 gruppering 1
14882 grupperingar 4
14883 grupperna 42
14884 gruppernas 1
14885 gruppers 5
14886 gruppkollega 1
14887 gruppkolleger 1
14888 gruppnivå 1
14889 gruppnivåer 2
14890 gruppnivån 2
14891 gruppordförande 1
14892 gruppordförandekommittén 1
14893 grupps 16
14894 grupptillhörighet 2
14895 gruppundantaget 1
14896 gruppvis 1
14897 gruva 2
14898 gruvan 1
14899 gruvbolaget 1
14900 gruvbolagets 1
14901 gruvbrytningen 1
14902 gruvbrytningens 1
14903 gruvbrytningsföretag 1
14904 gruvjobbarpub 1
14905 gruvnäringen 1
14906 gruvor 2
14907 grym 2
14908 grymhet 1
14909 grymt 5
14910 grymta 1
14911 grytor 1
14912 grytorna 1
14913 gräddtårtan 1
14914 gräl 4
14915 grälade 2
14916 grälar 1
14917 grämelse 1
14918 gränd 1
14919 gränden 2
14920 gräns 8
14921 gränsar 4
14922 gränsdragning 1
14923 gränsen 12
14924 gränser 54
14925 gränserna 38
14926 gränsfrågan 3
14927 gränskonflikter 1
14928 gränskontroll 3
14929 gränskontroller 2
14930 gränskontrollerna 1
14931 gränskontrollorganet 1
14932 gränskontrollsystemet 1
14933 gränslandet 1
14934 gränslinjen 1
14935 gränslöst 2
14936 gränsområde 2
14937 gränsområden 2
14938 gränsområdena 4
14939 gränsområdenas 1
14940 gränsprocesserna 1
14941 gränsregioner 2
14942 gränsregionerna 2
14943 gränsregionernas 1
14944 gränssmugglingen 1
14945 gränssnitt 1
14946 gränstrakterna 2
14947 gränsvärde 1
14948 gränsvärdena 1
14949 gränsövergripande 1
14950 gränsövergångsnivå 1
14951 gränsöverskridande 54
14952 gräset 3
14953 gräsligas 1
14954 gräslighet 1
14955 gräsligt 1
14956 gräsmatta 1
14957 gräsmattan 3
14958 gräsrotsgrupper 1
14959 gräsrotsnivå 1
14960 grässkjul 1
14961 grät 2
14962 gräver 2
14963 grävt 1
14964 grå 5
14965 grå- 1
14966 grådaskighet 1
14967 grånad 1
14968 gråt 2
14969 gråta 2
14970 grått 2
14971 gråvita 1
14972 gråzon 2
14973 grödor 1
14974 grön 12
14975 gröna 51
14976 grönare 1
14977 grönas 3
14978 grönbok 1
14979 grönböcker 1
14980 grönska 2
14981 grönskande 1
14982 grönt 3
14983 gröt 1
14984 grövsta 2
14985 gubbe 1
14986 gubben 4
14987 gud 3
14988 gudabild 1
14989 gudinna 1
14990 guds 3
14991 gudskelov 1
14992 gul 2
14993 gula 2
14994 gulag 1
14995 gulblekt 1
14996 gulbruna 1
14997 guld 4
14998 guldbokstäver 1
14999 gulden 1
15000 guldet 2
15001 guldgruva 1
15002 guldhöna 1
15003 guldringar 1
15004 gullegrisar 1
15005 gult 3
15006 gummidocka 1
15007 gummiparagraf 1
15008 gummistämpel 1
15009 gummistövlar 1
15010 gunga 1
15011 gungade 1
15012 gungades 1
15013 gungande 1
15014 gungar 1
15015 guvenörskap 1
15016 guvernör 2
15017 guvernören 1
15018 guvernörens 1
15019 gyllene 4
15020 gym 1
15021 gymnasiet 1
15022 gymnasium 1
15023 gynna 15
15024 gynnade 6
15025 gynnar 10
15026 gynnas 1
15027 gynnsam 4
15028 gynnsamma 7
15029 gynnsamt 1
15030 gyroskop 1
15031 gyttjemark 1
15032 gyttjig 1
15033 gyttjiga 1
15034 gäck 1
15035 gäldenärens 1
15036 gälla 47
15037 gällande 61
15038 gällde 24
15039 gäller 1022
15040 gällt 5
15041 gäng 2
15042 gängse 1
15043 gärna 122
15044 gärning 3
15045 gärningar 5
15046 gärningsmannen 1
15047 gärningsmän 2
15048 gäspa 1
15049 gäspade 1
15050 gäss 1
15051 gäst 4
15052 gäster 1
15053 gästerna 1
15054 gästfrihet 1
15055 gästhyddan 1
15056 gästrummet 1
15057 gå 238
15058 gång 244
15059 gångarna 3
15060 gången 81
15061 gånger 85
15062 gångna 8
15063 gångs 5
15064 går 310
15065 gård 1
15066 gårdagens 9
15067 gårdar 1
15068 gården 3
15069 gås 2
15070 gåsmarsch 1
15071 gåspenna 1
15072 gåta 4
15073 gåtan 1
15074 gåtfulla 1
15075 gåtfullt 2
15076 gått 61
15077 gåva 1
15078 göda 1
15079 gödsel 1
15080 gödseln 1
15081 gömda 1
15082 gömde 1
15083 gömma 2
15084 gömmas 1
15085 gömmer 5
15086 gömställe 1
15087 gömts 1
15088 gör 387
15089 göra 795
15090 göras 69
15091 görs 47
15092 ha 610
15093 habitat- 1
15094 habitatdirektiv 1
15095 habitatdirektivet 2
15096 hack 1
15097 hackande 1
15098 hade 691
15099 haft 88
15100 hajade 1
15101 hakat 1
15102 halka 1
15103 halkar 1
15104 hallen 4
15105 halm 2
15106 halogenerade 1
15107 hals 4
15108 halsar 1
15109 halsarna 1
15110 halsband 1
15111 halsbrytande 1
15112 halsduk 1
15113 halsen 5
15114 halt 2
15115 halta 1
15116 halte 1
15117 halv 12
15118 halva 10
15119 halvan 1
15120 halvdunklet 1
15121 halverades 1
15122 halverats 1
15123 halveringen 1
15124 halvhjärtade 1
15125 halvhjärtat 1
15126 halvideologiska 1
15127 halvkloten 1
15128 halvklädda 1
15129 halvmiljon 1
15130 halvoffentliga 1
15131 halvsovit 1
15132 halvt 6
15133 halvtidsbedömningen 1
15134 halvtimme 5
15135 halvvuxen 1
15136 halvvägs 6
15137 halvår 1
15138 halvåret 3
15139 halvårsskifte 1
15140 halvårsskiftet 2
15141 halvö 2
15142 halvön 2
15143 hamburgare 2
15144 hammare 2
15145 hamn 22
15146 hamna 7
15147 hamnade 3
15148 hamnanläggningen 1
15149 hamnar 47
15150 hamnarna 20
15151 hamnarnas 1
15152 hamnat 9
15153 hamnavgiften 2
15154 hamnavgifter 3
15155 hamnavgifterna 2
15156 hamnbestämmelser 1
15157 hamnen 19
15158 hamninspektioner 1
15159 hamnkategorier 1
15160 hamnkontroll 1
15161 hamnkontrollen 1
15162 hamnmyndigheterna 2
15163 hamnstaten 1
15164 hamra 1
15165 han 971
15166 hand 140
15167 handbagaget 1
15168 handdukar 1
15169 handel 36
15170 handeln 21
15171 handelns 1
15172 handels- 7
15173 handelsaspekter 1
15174 handelsavtal 9
15175 handelsavtalen 3
15176 handelsavtalet 6
15177 handelsavtalets 1
15178 handelsbalans 1
15179 handelsblockad 1
15180 handelsbolaget 1
15181 handelsfartyg 1
15182 handelsflotta 2
15183 handelsfrågor 3
15184 handelsförbindelser 1
15185 handelsförbindelserna 1
15186 handelsförhandlingar 1
15187 handelsförhandlingarna 1
15188 handelsförmåner 2
15189 handelsglobaliseringen 1
15190 handelshinder 2
15191 handelsintresseaspekten 1
15192 handelsintressen 1
15193 handelskrig 2
15194 handelslogik 1
15195 handelsmässiga 2
15196 handelsmässigt 1
15197 handelsområdet 1
15198 handelsplats 1
15199 handelsplatsen 1
15200 handelsplatser 1
15201 handelspolitik 4
15202 handelspolitiken 2
15203 handelsreformerna 1
15204 handelsregler 1
15205 handelsreglerna 1
15206 handelsrelaterade 1
15207 handelsrunda 1
15208 handelsrätt 2
15209 handelsrätten 1
15210 handelssamarbete 2
15211 handelssanktioner 1
15212 handelssektorn 1
15213 handelssidan 1
15214 handelssjöfart 1
15215 handelssjöfarten 1
15216 handelsstation 1
15217 handelstvisterna 1
15218 handelsuppgörelser 1
15219 handelsutbyte 4
15220 handelsutbyten 1
15221 handelsutbytespolitik 1
15222 handelsutbytet 3
15223 handelsutveckling 1
15224 handelsvara 4
15225 handelsystem 1
15226 handen 30
15227 handfast 1
15228 handfatet 1
15229 handflata 1
15230 handflatan 1
15231 handflator 1
15232 handfull 4
15233 handha 1
15234 handicap 1
15235 handikapp 8
15236 handikappade 9
15237 handikappades 4
15238 handla 20
15239 handlade 13
15240 handlande 5
15241 handlar 288
15242 handlare 1
15243 handlarna 1
15244 handlas 1
15245 handlat 3
15246 handling 34
15247 handlingar 41
15248 handlingarna 5
15249 handlingen 1
15250 handlingens 1
15251 handlingsalternativ 1
15252 handlingsansvar 1
15253 handlingsfrihet 1
15254 handlingsförlamning 1
15255 handlingsförmåga 3
15256 handlingsförmågan 1
15257 handlingskraft 4
15258 handlingskraftig 1
15259 handlingskraftiga 2
15260 handlingskraftigt 1
15261 handlingslinjer 3
15262 handlingsplan 14
15263 handlingsplanen 4
15264 handlingsplaner 8
15265 handlingsplanernas 1
15266 handlingsprogram 11
15267 handlingsramen 1
15268 handlingssätt 5
15269 handlingssätten 1
15270 handlingssättet 2
15271 handlingsutrymme 5
15272 handläggning 2
15273 handläggningen 2
15274 hands 2
15275 handskarna 1
15276 handskas 13
15277 handske 1
15278 handtaget 1
15279 handuppräckning 2
15280 handvändning 1
15281 handväska 1
15282 handväskan 1
15283 hankar 1
15284 hans 289
15285 hantera 40
15286 hanterande 1
15287 hanterandet 1
15288 hanterar 6
15289 hanteras 15
15290 hantering 22
15291 hanteringen 10
15292 hantlangare 1
15293 hantverk 2
15294 hantverkare 2
15295 hantverkarnas 1
15296 hantverksmässiga 2
15297 happy 1
15298 har 5034
15299 haranger 1
15300 haren 1
15301 harmoni 4
15302 harmoniera 1
15303 harmonisera 10
15304 harmoniserad 1
15305 harmoniserade 4
15306 harmoniserar 1
15307 harmoniseras 2
15308 harmoniserat 3
15309 harmoniserats 2
15310 harmonisering 40
15311 harmoniseringen 4
15312 harmoniseringsbegrepp 1
15313 harmonisk 10
15314 harmoniskt 1
15315 harpa 1
15316 hasande 2
15317 hasch 1
15318 hast 2
15319 hastigast 1
15320 hastighet 6
15321 hastigheten 2
15322 hastigheter 2
15323 hastigt 7
15324 hat 2
15325 hatade 1
15326 hatar 1
15327 hatet 3
15328 hatisk 1
15329 hatt 2
15330 hattar 3
15331 hattarna 1
15332 hatten 2
15333 hav 22
15334 havande 1
15335 have 1
15336 have-nots 2
15337 haven 12
15338 havens 2
15339 havererade 1
15340 haveri 5
15341 haveriet 1
15342 haves 2
15343 havet 64
15344 havets 9
15345 havs 23
15346 havs- 1
15347 havsbotten 1
15348 havsdimension 1
15349 havsdäggdjur 1
15350 havsfiske 1
15351 havsforskningsrådet 1
15352 havsföroreningar 2
15353 havsgränsen 1
15354 havsgränser 4
15355 havsgränserna 2
15356 havsinriktning 1
15357 havslivet 1
15358 havsmiljö 4
15359 havsmiljöer 1
15360 havsmiljön 8
15361 havsmiljöns 1
15362 havsnära 1
15363 havsområden 5
15364 havsområdena 1
15365 havsområdenas 1
15366 havsområdet 2
15367 havspolitik 1
15368 havsprodukternas 1
15369 havssköldpaddor 1
15370 havsströmmarna 1
15371 havsvattnet 2
15372 headline 2
15373 hearingen 1
15374 hebreiska 1
15375 heder 2
15376 hederliga 1
15377 hedersamt 1
15378 hederskompani 1
15379 hedersläktaren 1
15380 hedersmedlem 1
15381 hedervärt 2
15382 hedga 2
15383 hedniska 1
15384 hedra 5
15385 hedrade 2
15386 hedrande 1
15387 hedrar 1
15388 hejda 2
15389 hejdade 2
15390 hejdas 3
15391 hejdat 1
15392 hejdlösa 1
15393 hektar 3
15394 hektiska 1
15395 hektometer3 2
15396 hektona 1
15397 hel 42
15398 hela 415
15399 helgar 1
15400 helgdag 1
15401 helgdagar 1
15402 helgedom 1
15403 helgen 2
15404 helgjutna 1
15405 helgon 1
15406 helhet 57
15407 helheten 1
15408 helhetlig 1
15409 helhetsbalansen 1
15410 helhetsbild 1
15411 helhetskoncept 1
15412 helhetslösning 1
15413 helhetspolitik 1
15414 helhetssyn 1
15415 helhetssynen 1
15416 helhjärtad 1
15417 helhjärtade 1
15418 helhjärtat 10
15419 helig 1
15420 heliga 4
15421 helikopter 2
15422 helikoptern 1
15423 helikoptrar 7
15424 helikoptrarna 1
15425 heller 134
15426 hellre 14
15427 hellånga 1
15428 helsike 1
15429 helst 125
15430 helt 408
15431 heltidsanställning 1
15432 heltidsjobb 1
15433 heltäckande 8
15434 heltäckningsmattor 1
15435 helvete 2
15436 hem 47
15437 hemarbetet 1
15438 hembygd 1
15439 hemfalla 1
15440 hemförde 1
15441 hemifrån 1
15442 hemkommun 1
15443 hemkänsla 1
15444 hemkära 1
15445 hemland 14
15446 hemlandet 2
15447 hemlig 3
15448 hemliga 7
15449 hemlighet 4
15450 hemligheten 2
15451 hemligheter 3
15452 hemligheterna 1
15453 hemlighetsfulla 1
15454 hemlighetsfullt 3
15455 hemlighålla 2
15456 hemligt 1
15457 hemländer 2
15458 hemläxor 1
15459 hemlösa 7
15460 hemlöshet 3
15461 hemma 20
15462 hemmabasen 1
15463 hemmagjorda 1
15464 hemmamarknad 2
15465 hemmamarknader 2
15466 hemmaplan 1
15467 hemmasittare 1
15468 hemmet 5
15469 hemmets 1
15470 hemort 1
15471 hemregion 2
15472 hemsida 2
15473 hemsk 2
15474 hemska 6
15475 hemskaste 1
15476 hemskickad 1
15477 hemskt 1
15478 hemstad 1
15479 hemställer 1
15480 hemsökelser 1
15481 hemsökt 1
15482 hemvist 2
15483 hemväg 1
15484 henne 71
15485 hennes 84
15486 herodiska 1
15487 heroisk 1
15488 herr 490
15489 herrar 91
15490 herrarna 2
15491 herravälde 2
15492 herraväldet 1
15493 herrelösa 1
15494 herresäte 1
15495 herrgård 1
15496 herrtidningar 1
15497 hertigen 1
15498 hes 2
15499 het 3
15500 heta 6
15501 heter 13
15502 heterogena 1
15503 hets 2
15504 hetsen 1
15505 hett 6
15506 hetta 2
15507 hettan 3
15508 hette 6
15509 hexavalent 1
15510 hierarki 1
15511 hierarkin 2
15512 hierarkisering 1
15513 hierarkisk 1
15514 hierarkiska 1
15515 high 3
15516 himlen 6
15517 himmel 5
15518 himmelsskriande 1
15519 hinder 56
15520 hindra 17
15521 hindrade 3
15522 hindrades 1
15523 hindrar 28
15524 hindras 5
15525 hindrat 1
15526 hindrats 1
15527 hindren 3
15528 hindret 1
15529 hinduisk 1
15530 hink 1
15531 hinna 3
15532 hinner 1
15533 hisnande 1
15534 hissade 1
15535 hissen 1
15536 historia 42
15537 historien 15
15538 historiens 3
15539 historier 6
15540 historieskrivningen 1
15541 historik 1
15542 historiker 1
15543 historikern 1
15544 historisk 14
15545 historiska 20
15546 historiskt 12
15547 hit 35
15548 hitintills 1
15549 hitta 52
15550 hittade 6
15551 hittades 1
15552 hittar 12
15553 hittat 5
15554 hittats 1
15555 hittills 98
15556 hittillsvarande 6
15557 hiv-smitta 1
15558 hiv-smittade 1
15559 hivade 1
15560 hjord 2
15561 hjorden 1
15562 hjul 2
15563 hjulen 2
15564 hjulet 1
15565 hjulspår 1
15566 hjälm 1
15567 hjälp 165
15568 hjälpa 101
15569 hjälpande 3
15570 hjälpbehov 1
15571 hjälpen 11
15572 hjälper 12
15573 hjälpfunktion 1
15574 hjälpinsatsen 1
15575 hjälpinsatser 3
15576 hjälpkonstruktioner 1
15577 hjälplösa 2
15578 hjälpmedel 2
15579 hjälporganisationer 1
15580 hjälpprogram 1
15581 hjälpt 3
15582 hjälpta 1
15583 hjälpte 4
15584 hjälptjänster 1
15585 hjälpvilliga 1
15586 hjältar 1
15587 hjälten 1
15588 hjärna 1
15589 hjärnkapacitet 1
15590 hjärnor 2
15591 hjärnorna 1
15592 hjärta 7
15593 hjärtan 2
15594 hjärtans 3
15595 hjärtat 15
15596 hjärtliga 2
15597 hjärtligt 19
15598 hjärtpunkt 1
15599 hjässa 2
15600 hoande 1
15601 hobby 2
15602 hobbybilar 1
15603 hoc-direktiv 1
15604 hoc-transporter 1
15605 hojtade 1
15606 holländsk 1
15607 holländska 2
15608 home 1
15609 homofobin 1
15610 homogen 1
15611 homogena 1
15612 homogent 4
15613 homosexuell 1
15614 homosexuella 1
15615 hon 238
15616 honnör 1
15617 honom 243
15618 hop 1
15619 hopas 1
15620 hope 1
15621 hopfällbart 1
15622 hopkok 1
15623 hopp 19
15624 hoppa 2
15625 hoppade 1
15626 hoppades 7
15627 hoppar 1
15628 hoppas 284
15629 hoppats 1
15630 hoppet 5
15631 hoppfullhet 1
15632 hoppingivande 3
15633 hopplös 1
15634 hopplöst 6
15635 hora 1
15636 hord 1
15637 horderna 1
15638 horisont 1
15639 horisontala 2
15640 horisontella 3
15641 horisontellt 3
15642 horisonten 3
15643 hormonbehandlat 1
15644 hormonstörande 2
15645 horn 2
15646 hornen 1
15647 hos 185
15648 hospice 1
15649 hostade 2
15650 hot 31
15651 hota 2
15652 hotad 4
15653 hotade 6
15654 hotades 3
15655 hotande 4
15656 hotar 25
15657 hotas 15
15658 hotat 2
15659 hotats 2
15660 hotbilden 1
15661 hotbilder 1
15662 hotell 1
15663 hotell- 1
15664 hotellen 1
15665 hotellet 2
15666 hotellets 1
15667 hotellägare 1
15668 hotelser 2
15669 hotet 10
15670 hotfull 1
15671 hotfulla 1
15672 hotfullt 1
15673 hud 1
15674 huden 1
15675 hudfärg 3
15676 hugg 3
15677 hugga 1
15678 huggas 1
15679 hukade 2
15680 huliganerna 1
15681 human 2
15682 humanism 1
15683 humanistiska 2
15684 humanitet 1
15685 humanitär 14
15686 humanitära 19
15687 humanitäras 2
15688 humanitärt 4
15689 humankapital 3
15690 humankapitalet 1
15691 humlen 1
15692 humor 1
15693 humör 2
15694 hund 3
15695 hundar 1
15696 hundbajs 1
15697 hunden 2
15698 hundra 9
15699 hundrade 1
15700 hundrafemtio 1
15701 hundraprocentig 2
15702 hundraprocentigt 1
15703 hundraser 1
15704 hundratal 1
15705 hundratals 12
15706 hundratusentals 12
15707 hundskall 1
15708 hunger 1
15709 hungersnöd 2
15710 hungrig 3
15711 hunnit 4
15712 hur 537
15713 hurdan 2
15714 huruvida 27
15715 hus 26
15716 husalf 2
15717 husalfer 1
15718 husarrest 1
15719 husbonde 1
15720 husdjur 1
15721 husen 2
15722 huset 19
15723 husets 2
15724 hushåll 4
15725 hushålla 1
15726 hushållen 1
15727 hushållning 2
15728 hushålls- 1
15729 hushållsvatten 1
15730 hushållsändamål 1
15731 husligt 1
15732 husrum 1
15733 hustak 1
15734 hustru 15
15735 hustrun 3
15736 hustruns 1
15737 husövertaganden 1
15738 huva 1
15739 huvan 1
15740 huvud 35
15741 huvudaktiviteter 1
15742 huvudaktör 1
15743 huvudangelägenheter 1
15744 huvudansvaret 5
15745 huvudargument 1
15746 huvudbeståndsdelar 1
15747 huvudbudskap 2
15748 huvudbyggnad 1
15749 huvuddel 1
15750 huvuddelen 1
15751 huvuddrag 1
15752 huvuddragen 3
15753 huvuden 3
15754 huvudena 1
15755 huvudet 17
15756 huvudfinansieringen 1
15757 huvudfråga 4
15758 huvudfrågan 1
15759 huvudförslagen 1
15760 huvudinriktning 1
15761 huvudinriktningar 1
15762 huvudkontor 3
15763 huvudkravet 1
15764 huvudlinjerna 2
15765 huvudmål 3
15766 huvudpersonerna 1
15767 huvudprincip 1
15768 huvudpunkter 1
15769 huvudrekommendationer 1
15770 huvudroll 3
15771 huvudrollsinnehavarna 1
15772 huvudrubriker 1
15773 huvudsak 18
15774 huvudsaken 2
15775 huvudsakliga 15
15776 huvudsaklige 1
15777 huvudsakligen 30
15778 huvudskälet 1
15779 huvudstad 4
15780 huvudstaden 1
15781 huvudstadens 1
15782 huvudstäder 2
15783 huvudstäderna 3
15784 huvudsyfte 1
15785 huvudsyften 1
15786 huvudsyftet 1
15787 huvudtaget 1
15788 huvuduppgift 1
15789 huvuduppgifter 1
15790 huvudvärk 2
15791 hy 5
15792 hybridbetänkande 1
15793 hycklade 1
15794 hycklande 4
15795 hyckleri 8
15796 hyckleriet 2
15797 hyddan 1
15798 hyddor 2
15799 hydrauliska 1
15800 hydrogeologiskt 1
15801 hydrologiska 1
15802 hygglig 1
15803 hygien 3
15804 hygienens 1
15805 hygieniska 1
15806 hylla 5
15807 hyllade 1
15808 hyllan 1
15809 hyllandet 1
15810 hyllar 1
15811 hyllas 1
15812 hyllning 2
15813 hylsa 1
15814 hypereffektiva 1
15815 hypnotiserade 1
15816 hypotes 1
15817 hypotesen 1
15818 hypoteser 1
15819 hypotetiska 1
15820 hypotetiskt 2
15821 hyr 1
15822 hyrd 1
15823 hyreshus 1
15824 hysa 7
15825 hyser 10
15826 hyste 1
15827 hysterin 1
15828 hytt 1
15829 hytten 2
15830 häcken 5
15831 hädanefter 2
15832 hädelser 2
15833 häftiga 4
15834 häftigt 2
15835 hägn 1
15836 häktade 1
15837 häktningen 1
15838 häktningsorder 1
15839 häl 1
15840 häleri 1
15841 hälft 2
15842 hälften 17
15843 hällde 1
15844 hälsa 50
15845 hälsade 6
15846 hälsades 1
15847 hälsan 8
15848 hälsar 9
15849 hälsning 1
15850 hälsningar 2
15851 hälsningen 1
15852 hälso- 6
15853 hälsoaspekten 1
15854 hälsobehoven 1
15855 hälsobringande 1
15856 hälsoeffekter 1
15857 hälsoeffekterna 1
15858 hälsofrämjande 1
15859 hälsofrågor 3
15860 hälsoområden 1
15861 hälsoproblem 1
15862 hälsoproblemen 1
15863 hälsorelaterade 1
15864 hälsorisker 1
15865 hälsosam 2
15866 hälsosamma 1
15867 hälsosektorn 3
15868 hälsosituationen 1
15869 hälsoskydd 3
15870 hälsoskyddet 1
15871 hälsosystemet 1
15872 hälsotillstånd 3
15873 hälsotjänster 1
15874 hälsovådliga 1
15875 hälsovård 13
15876 hälsovården 3
15877 hälsovårdsanordningar 1
15878 hälsovårdsdepartement 1
15879 hälsovårdsinrättningar 2
15880 hälsovårdsinspektören 1
15881 hälsovårdskostnader 1
15882 hälsovårdsområdet 1
15883 hälsovårdssystem 2
15884 hälsovårdssystemet 3
15885 hämma 1
15886 hämmar 2
15887 hämmas 1
15888 hämnande 1
15889 hämnas 2
15890 hämnd 2
15891 hämndbegär 1
15892 hämndlystnad 1
15893 hämningslös 1
15894 hämta 8
15895 hämtad 1
15896 hämtade 2
15897 hämtar 2
15898 hämtas 4
15899 hämtat 2
15900 hämtning 1
15901 hända 31
15902 hände 31
15903 händelse 30
15904 händelseförloppet 1
15905 händelselös 1
15906 händelsemönster 1
15907 händelsen 6
15908 händelsens 1
15909 händelser 37
15910 händelserikt 1
15911 händelserna 17
15912 händelseutveckling 1
15913 händelseutvecklingen 1
15914 händelsevis 2
15915 händer 54
15916 händerna 22
15917 händigt 1
15918 hänför 2
15919 hänförde 1
15920 hänga 5
15921 hängande 4
15922 hängbro 1
15923 hängde 14
15924 hänge 1
15925 hänger 28
15926 hängett 1
15927 hängivelse 1
15928 hängivenhet 1
15929 hänglås 1
15930 hängning 1
15931 hängslen 1
15932 hänseende 15
15933 hänseenden 4
15934 hänseendet 4
15935 hänskjuta 1
15936 hänsyn 199
15937 hänsynen 5
15938 hänsynsfull 1
15939 hänsynstaganden 3
15940 hänsynstagandet 3
15941 hänt 26
15942 hänvisa 20
15943 hänvisad 1
15944 hänvisade 18
15945 hänvisades 2
15946 hänvisar 22
15947 hänvisas 5
15948 hänvisat 6
15949 hänvisats 3
15950 hänvisning 22
15951 hänvisningar 8
15952 hänvisningarna 1
15953 hänvisningen 8
15954 häpen 1
15955 häpnad 3
15956 häpnadsväckande 1
15957 häpnar 1
15958 här 1129
15959 härden 1
15960 härefter 1
15961 häri 1
15962 härifrån 3
15963 härigenom 4
15964 härjade 2
15965 härledas 2
15966 härliga 1
15967 härligaste 1
15968 härligt 1
15969 härmade 2
15970 härmed 11
15971 häromdagen 1
15972 härrör 19
15973 härs 1
15974 härskar 1
15975 härskare 2
15976 härskarinnan 1
15977 härskarna 1
15978 härskaror 1
15979 härstammar 7
15980 härtill 1
15981 härutöver 1
15982 härva 1
15983 härvidlag 1
15984 häst 5
15985 hästar 2
15986 hästen 4
15987 hästliknande 1
15988 hästskor 1
15989 häva 5
15990 hävas 3
15991 hävda 18
15992 hävdade 8
15993 hävdar 22
15994 hävdas 1
15995 hävdat 7
15996 hävdvunna 1
15997 häver 2
15998 hävning 1
15999 hävstången 1
16000 hävts 1
16001 häxa 3
16002 häxan 1
16003 häxkonst 1
16004 häxkonster 1
16005 häxor 1
16006 hågen 1
16007 håglöst 1
16008 hål 5
16009 håla 1
16010 håll 46
16011 hålla 96
16012 hållas 14
16013 hållbar 85
16014 hållbara 15
16015 hållbarhet 5
16016 hållbart 18
16017 hållen 2
16018 håller 186
16019 hållet 38
16020 hållit 17
16021 hållits 3
16022 hållna 2
16023 hållning 24
16024 hållningen 2
16025 hållplats 1
16026 hålls 13
16027 hålor 1
16028 hån 2
16029 hånade 1
16030 hånar 1
16031 hånflinande 1
16032 hånfull 1
16033 hår 17
16034 hård 13
16035 hårda 15
16036 hårdare 5
16037 hårdast 4
16038 hårdhandskarna 1
16039 hårdingar 1
16040 hårdingen 1
16041 hårdnackade 1
16042 hårdnackat 2
16043 håret 10
16044 hårfina 1
16045 hårklyverier 1
16046 hårnät 1
16047 hårnål 1
16048 hårnålar 1
16049 hårnålen 1
16050 hårstrå 2
16051 hårt 46
16052 hårtestar 1
16053 håvar 1
16054 höft 1
16055 höfterna 1
16056 hög 104
16057 höga 60
16058 högaktar 1
16059 högaktuellt 1
16060 högar 1
16061 höge 34
16062 höger 12
16063 högerextremismen 1
16064 högerextremismens 1
16065 högerextremistiska 3
16066 högerhanden 1
16067 högerkanten 1
16068 högerkvinnor 1
16069 högerledamöters 1
16070 högermajoritet 1
16071 högern 5
16072 högerns 4
16073 högerpopulists 1
16074 högervridning 1
16075 högg 1
16076 höghastighetståg 1
16077 höginkomstländer 1
16078 höginkomsttagare 1
16079 högkonjunktur 1
16080 högkostnadsområden 1
16081 högkvalitativ 2
16082 högkvalitativa 1
16083 högkvarter 1
16084 högljudd 1
16085 högljudda 1
16086 högljutt 2
16087 högländerna 2
16088 högnivågrupp 3
16089 högnivågruppen 6
16090 högprestationstjänst 1
16091 högpresterande 1
16092 högra 1
16093 högre 77
16094 högrest 1
16095 högriskfonder 1
16096 högriskprodukter 1
16097 högröda 1
16098 högrörliga 1
16099 högskolor 1
16100 högst 37
16101 högsta 38
16102 högste 1
16103 högstämda 1
16104 högt 38
16105 högteknologiska 2
16106 högtidliga 1
16107 högtidligen 1
16108 högtidligheten 1
16109 högtidlighålla 1
16110 högtidligt 8
16111 högtravande 2
16112 höja 15
16113 höjas 5
16114 höjd 8
16115 höjda 2
16116 höjde 2
16117 höjden 1
16118 höjderna 1
16119 höjdpunkt 2
16120 höjdpunkten 1
16121 höjer 3
16122 höjning 7
16123 höjningar 1
16124 höjningen 3
16125 höjs 2
16126 höjt 1
16127 höjts 1
16128 hölje 1
16129 höljs 1
16130 höll 37
16131 hölls 5
16132 höna 1
16133 hönor 1
16134 hör 90
16135 höra 70
16136 hörande 1
16137 höras 5
16138 hörbar 1
16139 hörbart 1
16140 hörd 4
16141 hörda 1
16142 hörde 33
16143 hördes 10
16144 hörn 4
16145 hörnen 2
16146 hörnet 4
16147 hörnsten 2
16148 hörnstenen 1
16149 hörsammar 1
16150 hörsammats 2
16151 hört 74
16152 hörts 3
16153 höst 2
16154 höstack 1
16155 höstas 2
16156 hösten 3
16157 hövlig 1
16158 hövlighet 1
16159 i 12516
16160 i- 1
16161 iaktta 10
16162 iakttagande 4
16163 iakttagelse 1
16164 iakttagelser 4
16165 iakttagelserna 1
16166 iakttagit 1
16167 iakttar 2
16168 iakttas 6
16169 iakttog 3
16170 ianspråktagandet 1
16171 iberiska 1
16172 ibland 59
16173 icke 41
16174 icke- 1
16175 icke-albaner 1
16176 icke-albanska 3
16177 icke-avvisning 1
16178 icke-bergsregioner 1
16179 icke-budgetisering 1
16180 icke-danska 1
16181 icke-diskriminerande 1
16182 icke-diskriminering 3
16183 icke-dokument 1
16184 icke-européer- 1
16185 icke-fossil 1
16186 icke-handikappade 1
16187 icke-harmoniserade 3
16188 icke-inblandning 1
16189 icke-införlivande 1
16190 icke-insatta 1
16191 icke-intervention 1
16192 icke-interventionsmotionen 1
16193 icke-kommersiella 1
16194 icke-kvalificerade 1
16195 icke-lönerelaterade 1
16196 icke-medborgare 1
16197 icke-medlemsstater 1
16198 icke-metalldelar 1
16199 icke-militära 1
16200 icke-rasistiskt 1
16201 icke-regeringssektorns 1
16202 icke-självvalda 1
16203 icke-spridningsavtalet 3
16204 icke-statlig 1
16205 icke-statliga 40
16206 icke-statligt 1
16207 icke-tariffiära 1
16208 icke-tillämpning 1
16209 icke-ömsesidiga 1
16210 ickenylonhud 1
16211 ickesjälsligt 1
16212 idag 12
16213 ideal 4
16214 ideala 2
16215 idealen 2
16216 idealet 2
16217 idealiserat 1
16218 idealisk 1
16219 idealiska 1
16220 idealiskt 1
16221 idealism 2
16222 idealistiskt 1
16223 ideella 2
16224 idel 1
16225 ideligen 2
16226 identifiera 13
16227 identifierade 4
16228 identifierades 1
16229 identifierar 5
16230 identifieras 4
16231 identifierat 6
16232 identifierats 1
16233 identifierbara 1
16234 identifiering 1
16235 identifieringen 1
16236 identifikation 1
16237 identisk 1
16238 identiska 1
16239 identiskt 1
16240 identitet 15
16241 identiteten 3
16242 identiteter 2
16243 identitetshandlingar 2
16244 ideolog 1
16245 ideologi 4
16246 ideologisk 2
16247 ideologiska 7
16248 ideologiskt 2
16249 idiosynkrasi 1
16250 idiot 3
16251 idiotiska 1
16252 idrott 5
16253 idrottssammanhang 1
16254 idyllisk 1
16255 idé 26
16256 idéer 34
16257 idéerna 1
16258 idén 32
16259 ifall 7
16260 ifråga 3
16261 ifrågasatt 1
16262 ifrågasatte 1
16263 ifrågasattes 2
16264 ifrågasatts 1
16265 ifrågasätta 13
16266 ifrågasättande 3
16267 ifrågasättanden 1
16268 ifrågasättandet 1
16269 ifrågasättas 4
16270 ifrågasätter 12
16271 ifrågasätts 6
16272 ifrågavarande 4
16273 ifrån 74
16274 iförd 4
16275 igelkott 1
16276 igen 127
16277 igenkännande 3
16278 igenom 67
16279 igenom- 1
16280 igenspikade 1
16281 ignorera 4
16282 ignorerade 2
16283 ignorerades 1
16284 ignoreras 3
16285 igång 29
16286 igångkörning 1
16287 igångsättandet 2
16288 ihjäl 1
16289 ihop 48
16290 ihärdighet 1
16291 ihåg 45
16292 ihåliga 1
16293 ihållande 8
16294 ikapp 1
16295 ikraftträdande 4
16296 ikraftträdandet 3
16297 il 1
16298 illa 16
16299 illaluktande 1
16300 illavarslande 2
16301 illegal 5
16302 illegala 12
16303 illegalt 5
16304 illojal 1
16305 illojala 2
16306 illusion 4
16307 illusionen 1
16308 illusioner 1
16309 illusionism 1
16310 illusionsfrie 1
16311 illusoriskt 1
16312 illustration 2
16313 illustrera 3
16314 illustrerade 1
16315 illustrerar 1
16316 illustreras 2
16317 illvilliga 1
16318 illvilligt 1
16319 ilska 3
16320 ilsken 1
16321 ilsket 3
16322 ilskna 2
16323 image 1
16324 imaginära 1
16325 imitationsprodukter 1
16326 imitera 1
16327 immaterialrätt 3
16328 immaterialrätten 3
16329 immaterialrättsliga 2
16330 immaterialrättsligt 2
16331 immateriella 5
16332 immigrantbefolkningen 1
16333 immigranter 3
16334 immigration 3
16335 immigrationen 1
16336 immigrationsblanketterna 1
16337 immigrationspolitiken 1
16338 immigrationsprocess 1
16339 immunitet 7
16340 immuniteten 5
16341 imperativ 2
16342 imperialisternas 1
16343 imperialistiska 1
16344 imperiebyggare 1
16345 implementation 1
16346 implementerade 2
16347 implementeringen 2
16348 implicit 1
16349 imponera 1
16350 imponerad 1
16351 imponerade 1
16352 imponerande 3
16353 impopulärt 1
16354 import 6
16355 importbegränsningarna 1
16356 importen 5
16357 importera 3
16358 importerad 3
16359 importerade 3
16360 importerar 1
16361 importeras 4
16362 importerats 1
16363 importförbudet 1
16364 importhinder 1
16365 importpolitik 2
16366 importrestriktioner 1
16367 importsystemet 1
16368 impossible 1
16369 improviserat 1
16370 impuls 3
16371 impulsen 1
16372 impulser 11
16373 impulsiv 1
16374 impunity 1
16375 in 400
16376 in- 1
16377 inaktiverat 1
16378 inaktivt 1
16379 inarbetats 1
16380 inbegripa 6
16381 inbegripande 1
16382 inbegripandet 1
16383 inbegripas 3
16384 inbegripen 1
16385 inbegriper 18
16386 inbegripet 20
16387 inbegripna 2
16388 inbegrips 2
16389 inbesparingar 1
16390 inbilla 2
16391 inbillad 1
16392 inbillade 1
16393 inbjuda 2
16394 inbjudan 2
16395 inbjudande 1
16396 inbjuden 2
16397 inbjuder 3
16398 inbjudit 1
16399 inbjudits 1
16400 inbjudna 2
16401 inbjudningar 1
16402 inbjöd 1
16403 inblandad 3
16404 inblandade 19
16405 inblandat 2
16406 inblandning 22
16407 inbringade 2
16408 inbringar 1
16409 inbyggd 2
16410 inbördes 21
16411 inbördeskrig 3
16412 inbördeskriget 2
16413 incident 1
16414 incitament 12
16415 incitamenten 1
16416 incitamentet 4
16417 indelade 2
16418 indelas 2
16419 indelat 1
16420 index 2
16421 indexering 1
16422 indexet 1
16423 indexfond 1
16424 indianer 1
16425 indianerna 2
16426 indianernas 1
16427 indianska 1
16428 indicier 2
16429 indignation 1
16430 indikation 1
16431 indikationer 1
16432 indikativt 1
16433 indikatorer 12
16434 indikatorn 1
16435 indirekt 15
16436 indirekta 6
16437 indiska 2
16438 individ 7
16439 individen 1
16440 individens 3
16441 individer 9
16442 individerna 1
16443 individers 1
16444 individs 1
16445 individualiserade 1
16446 individualisering 1
16447 individualism 2
16448 individualitet 1
16449 individuell 2
16450 individuella 14
16451 individuellt 2
16452 indonesisk 1
16453 indonesiska 1
16454 indonesiskt 1
16455 indraget 1
16456 indragning 1
16457 indränkt 1
16458 industri 16
16459 industri- 4
16460 industrial 1
16461 industrialiserade 2
16462 industrialiseringen 1
16463 industriell 2
16464 industriella 11
16465 industriellt 1
16466 industrier 7
16467 industrierna 1
16468 industriernas 1
16469 industrifrågor 6
16470 industriföretagen 1
16471 industriföroreningar 1
16472 industrigrupper 1
16473 industrikatastrofer 1
16474 industrikulturen 1
16475 industriliknande 1
16476 industrilobbyisten 1
16477 industriländerna 2
16478 industrimässor 1
16479 industrin 38
16480 industrins 4
16481 industripolitikerna 1
16482 industripolitisk 1
16483 industriprodukt 1
16484 industriprodukter 1
16485 industris 1
16486 industrisektorer 1
16487 industriverksamheten 1
16488 industriverksamheter 1
16489 indämda 1
16490 ineffektiv 2
16491 ineffektiva 4
16492 ineffektivitet 4
16493 ineffektivt 2
16494 infallsvinklar 1
16495 infallsvinklarna 1
16496 infann 1
16497 infantiliserande 1
16498 infekterade 2
16499 infektion 1
16500 infektionsnivåer 1
16501 infektionssjukdom 1
16502 infektiös 5
16503 infernaliska 2
16504 inferno 2
16505 infernos 1
16506 infiltrera 1
16507 infinitum 1
16508 infinner 1
16509 inflation 6
16510 inflationen 8
16511 inflationsbekämpning 1
16512 inflationsbekämpningen 1
16513 inflationstrycket 1
16514 influerad 1
16515 inflytande 23
16516 inflytelserika 1
16517 infogas 1
16518 information 145
16519 informationen 38
16520 informationer 1
16521 informations- 13
16522 informationsanalys 1
16523 informationsanalytiker 1
16524 informationsbrist 1
16525 informationsbudget 2
16526 informationsbärare 1
16527 informationscentrerna 1
16528 informationscentrum 1
16529 informationsekonomi 1
16530 informationsfattiga 1
16531 informationsflöde 1
16532 informationsfrihet 2
16533 informationsfrågan 1
16534 informationsinsamling 2
16535 informationskampanj 4
16536 informationskampanjen 2
16537 informationskampanjer 1
16538 informationskanal 1
16539 informationsmöte 1
16540 informationspolitik 1
16541 informationspolitiken 1
16542 informationsproblem 1
16543 informationsrika 1
16544 informationssamhälle 2
16545 informationssamhället 16
16546 informationssamhällets 1
16547 informationssystem 7
16548 informationsteknik 6
16549 informationstekniken 6
16550 informationsteknikmarknaderna 1
16551 informationsteknisk 1
16552 informationstekniska 2
16553 informationsteknologi 1
16554 informationsteknologin 4
16555 informationsutbyte 5
16556 informationsutbytet 4
16557 informationsvilja 1
16558 informationsåtgärder 2
16559 informationsöverföringens 1
16560 informella 7
16561 informellt 2
16562 informera 30
16563 informerad 3
16564 informerade 10
16565 informerades 2
16566 informerar 1
16567 informeras 6
16568 informerat 5
16569 informerats 3
16570 infrastruktur 21
16571 infrastrukturbestämmelser 1
16572 infrastrukturell 1
16573 infrastrukturella 1
16574 infrastrukturen 7
16575 infrastrukturens 2
16576 infrastrukturer 11
16577 infrastrukturerna 2
16578 infrastrukturnätet 1
16579 infrastrukturprogram 1
16580 infrastrukturprojekt 1
16581 infrastruktursatsningar 1
16582 infrastrukturutvecklingen 1
16583 infrastrukturåtgärder 1
16584 infria 1
16585 infriade 1
16586 infriades 1
16587 infrias 1
16588 infunnit 2
16589 infångad 1
16590 infödingarna 1
16591 inföll 1
16592 inför 279
16593 införa 94
16594 införande 8
16595 införandet 22
16596 införas 18
16597 införde 3
16598 infördes 5
16599 införliva 16
16600 införlivade 1
16601 införlivades 4
16602 införlivande 11
16603 införlivandet 9
16604 införlivar 3
16605 införlivas 15
16606 införlivat 1
16607 införlivats 5
16608 införs 9
16609 införsel 2
16610 införselrestriktioner 1
16611 införstådd 2
16612 införstådda 1
16613 infört 11
16614 införts 7
16615 inga 99
16616 ingalunda 6
16617 ingav 2
16618 ingavs 2
16619 inge 2
16620 ingen 214
16621 ingenjör 2
16622 ingenjörer 1
16623 ingenstans 4
16624 ingenting 85
16625 inger 6
16626 inget 90
16627 ingett 2
16628 ingick 3
16629 ingivit 8
16630 ingivits 3
16631 ingjuta 1
16632 ingrediens 1
16633 ingredienser 3
16634 ingrep 1
16635 ingrepp 9
16636 ingreppen 2
16637 ingress 1
16638 ingressen 1
16639 ingripa 20
16640 ingripande 13
16641 ingripanden 1
16642 ingripandet 1
16643 ingriper 3
16644 ingripit 4
16645 ingrott 1
16646 ingå 24
16647 ingående 14
16648 ingår 48
16649 ingått 8
16650 ingåtts 4
16651 inhemsk 1
16652 inhemska 11
16653 inhämta 2
16654 inhämtande 1
16655 inhämtar 1
16656 inhämtas 1
16657 inhämtat 1
16658 inifrån 4
16659 initiativ 161
16660 initiativandan 1
16661 initiativbetänkande 2
16662 initiativen 7
16663 initiativet 35
16664 initiativets 1
16665 initiativförmåga 1
16666 initiativkraft 2
16667 initiativrik 1
16668 initiativrikt 1
16669 initiativrätt 8
16670 initiativrätten 2
16671 initiativs 1
16672 initiativtagares 1
16673 initiera 1
16674 initierade 1
16675 initierades 1
16676 initierat 3
16677 injicerats 1
16678 inkapslade 2
16679 inkarnationen 2
16680 inkilade 1
16681 inkludera 11
16682 inkluderade 1
16683 inkluderades 1
16684 inkluderandet 1
16685 inkluderar 5
16686 inkluderas 5
16687 inkluderat 3
16688 inkluderats 1
16689 inklusive 47
16690 inkom 1
16691 inkompetens 3
16692 inkompetensen 1
16693 inkompetenta 1
16694 inkomst 7
16695 inkomst- 1
16696 inkomsten 2
16697 inkomster 17
16698 inkomsterna 3
16699 inkomstfördelning 1
16700 inkomstförluster 1
16701 inkomstkälla 4
16702 inkomstkällor 1
16703 inkomstskapande 1
16704 inkomststöd 1
16705 inkonsekvens 1
16706 inkonsekvenser 1
16707 inkonsekvenserna 1
16708 inkonsekvent 1
16709 inkorporera 1
16710 inkorrekta 1
16711 inkräkta 1
16712 inkubationsperiod 1
16713 inköp 3
16714 inköpsbesluten 1
16715 inköpslistor 2
16716 inköpslistorna 1
16717 inkörsport 1
16718 inlandet 1
16719 inlands- 1
16720 inlandsstaterna 1
16721 inleda 61
16722 inledande 7
16723 inledandet 2
16724 inledas 9
16725 inledde 9
16726 inleddes 11
16727 inleder 12
16728 inledning 1
16729 inledningen 10
16730 inledningsanförande 1
16731 inledningsfasen 1
16732 inledningsskedet 3
16733 inledningsvis 8
16734 inleds 12
16735 inlett 10
16736 inletts 20
16737 inlägg 42
16738 inlägga 1
16739 inläggen 4
16740 inlägget 2
16741 inlämnade 2
16742 inlämnades 2
16743 inlämnande 1
16744 inlämning 3
16745 inlämnings- 1
16746 inlämningsdatumen 1
16747 inlärningsproblem 1
16748 inlåsta 1
16749 inlåta 1
16750 inlåter 1
16751 inlöpande 1
16752 innan 124
16753 innandömen 2
16754 innanför 7
16755 inne 24
16756 inne-semantik 1
16757 innebar 8
16758 inneboende 3
16759 inneburit 3
16760 innebär 254
16761 innebära 59
16762 innebörd 4
16763 innebörden 12
16764 innefatta 1
16765 innefattade 1
16766 innefattande 1
16767 innefattar 12
16768 innefattas 8
16769 innehaft 1
16770 innehar 12
16771 innehas 2
16772 innehav 1
16773 innehavarna 1
16774 innehåll 30
16775 innehålla 16
16776 innehållande 2
16777 innehåller 97
16778 innehållet 51
16779 innehållit 2
16780 innehållsdeklaration 1
16781 innehållsindustrin 1
16782 innehållslig 1
16783 innehållsliga 3
16784 innehållsmässigt 2
16785 innehållsrika 2
16786 innehöll 9
16787 inneperiod 1
16788 innerfickan 1
16789 innerliga 3
16790 innerligt 3
16791 innerst 1
16792 innersta 2
16793 innerstad 1
16794 innersulor 1
16795 innevarande 3
16796 innevånare 2
16797 innovation 16
16798 innovationer 4
16799 innovationsföretag 1
16800 innovationspolitik 1
16801 innovationsprojekt 1
16802 innovativ 5
16803 innovativa 14
16804 innovativt 1
16805 innovatörer 1
16806 innovatörerna 1
16807 inofficiella 1
16808 inom 888
16809 inombords 1
16810 inomeuropeiska 1
16811 inomhustoalett 1
16812 inpränta 1
16813 inpräntat 1
16814 inpå 2
16815 inramad 1
16816 inramade 2
16817 inramning 2
16818 inre 201
16819 inresa 3
16820 inrikes 21
16821 inrikes- 3
16822 inrikesfrågor 2
16823 inrikesminister 1
16824 inrikesministeriet 1
16825 inrikesministern 3
16826 inrikesministrar 1
16827 inrikesministrarna 1
16828 inrikespolitik 3
16829 inrikespolitiska 3
16830 inrikta 14
16831 inriktad 10
16832 inriktade 5
16833 inriktar 5
16834 inriktas 5
16835 inriktat 5
16836 inriktning 32
16837 inriktningar 5
16838 inriktningen 10
16839 inrotad 1
16840 inryms 2
16841 inrätta 54
16842 inrättade 4
16843 inrättades 6
16844 inrättande 5
16845 inrättandet 21
16846 inrättar 6
16847 inrättas 13
16848 inrättat 3
16849 inrättats 5
16850 inrättningar 4
16851 inrättningarna 2
16852 inrådan 1
16853 insamlade 2
16854 insamlas 2
16855 insamling 19
16856 insamlingen 2
16857 insamlingsanläggning 1
16858 insamlingsmetoderna 1
16859 insats 35
16860 insatsen 3
16861 insatser 75
16862 insatserna 20
16863 insatsområden 1
16864 insatsområdena 1
16865 insatsstyrka 3
16866 insatsstyrkan 4
16867 insatt 1
16868 inse 32
16869 insegel 1
16870 insekter 2
16871 insektsmedel 1
16872 inser 41
16873 insett 3
16874 insikt 4
16875 insikten 4
16876 insikter 1
16877 insiktsfulla 1
16878 insistera 16
16879 insisterade 2
16880 insisterar 9
16881 inskickandet 1
16882 inskrida 1
16883 inskriven 2
16884 inskränka 6
16885 inskränkande 1
16886 inskränker 7
16887 inskränkning 3
16888 inskränkningar 4
16889 inskränkningarna 2
16890 inskränks 1
16891 inskränkte 1
16892 inskränkts 1
16893 inslag 11
16894 inslagen 3
16895 inslaget 2
16896 inslagna 2
16897 insläppningsknappen 1
16898 insolvens 4
16899 insolvensförfarande 1
16900 insolvensförfaranden 2
16901 inspekterades 1
16902 inspekteras 1
16903 inspektion 2
16904 inspektioner 4
16905 inspektionerna 1
16906 inspektionsmyndigheterna 1
16907 inspektionssystem 1
16908 inspektörer 5
16909 inspektörernas 1
16910 inspektörskår 1
16911 inspiration 1
16912 inspirationskällor 1
16913 inspiratörer 1
16914 inspirerad 1
16915 inspirerande 1
16916 inspireras 1
16917 inspirerat 1
16918 inspirerats 1
16919 inspärrade 1
16920 instabil 3
16921 instabila 1
16922 instabilitet 3
16923 instabiliteten 1
16924 installationerna 1
16925 installationsalternativ 1
16926 installationssidan 1
16927 installera 4
16928 installerade 1
16929 installeras 4
16930 installerat 4
16931 installerats 2
16932 instans 5
16933 instanser 9
16934 instanserna 7
16935 insteg 1
16936 instifta 2
16937 instiftats 1
16938 instinkt 1
16939 instinkter 1
16940 instinktiva 1
16941 instituten 2
16942 institution 28
16943 institutionell 9
16944 institutionella 32
16945 institutionellt 3
16946 institutionen 3
16947 institutionens 1
16948 institutioner 94
16949 institutionerna 76
16950 institutionernas 12
16951 institutioners 7
16952 institutionsansvariga 1
16953 institutionsprojekt 1
16954 institutionsreformen 1
16955 instruktioner 2
16956 instrument 110
16957 instrumentaliseras 1
16958 instrumentbrädan 1
16959 instrumenten 10
16960 instrumenterad 1
16961 instrumentet 15
16962 instrumentets 1
16963 instruments 2
16964 inställa 4
16965 inställd 9
16966 inställda 4
16967 inställer 3
16968 inställning 54
16969 inställningar 1
16970 inställningen 9
16971 inställsamma 1
16972 inställsamt 2
16973 inställt 2
16974 instämde 2
16975 instämma 13
16976 instämmande 4
16977 instämmer 41
16978 instängd 1
16979 instängda 2
16980 instängt 1
16981 insvept 1
16982 insyn 23
16983 insynen 3
16984 insynsskyddat 1
16985 insändare 1
16986 insättande 1
16987 insättningar 1
16988 insåg 8
16989 inta 14
16990 intagit 6
16991 intagits 1
16992 intakta 1
16993 intala 1
16994 intar 13
16995 intas 2
16996 inte 5114
16997 integration 26
16998 integrationen 20
16999 integrationens 2
17000 integrationsfaktor 1
17001 integrationsförfarande 1
17002 integrationsförmåga 1
17003 integrationsmekanismer 1
17004 integrationsmodellen 1
17005 integrationspolitik 3
17006 integrationsproblem 1
17007 integrationsprocess 2
17008 integrationsprocessen 5
17009 integrationsprogram 1
17010 integrationsstrategi 1
17011 integrationsåtgärderna 1
17012 integrera 19
17013 integrerad 14
17014 integrerade 4
17015 integrerades 1
17016 integrerandet 1
17017 integrerar 3
17018 integreras 13
17019 integrerat 5
17020 integrerats 1
17021 integrering 28
17022 integreringen 7
17023 integreringsarbetet 1
17024 integreringsprocesser 1
17025 integritet 6
17026 integriteten 1
17027 intellektuell 2
17028 intellektuella 6
17029 intellektuellt 3
17030 intelligens 1
17031 intelligensen 1
17032 intelligent 6
17033 intelligenta 2
17034 intensifiera 5
17035 intensifieras 1
17036 intensifieringen 1
17037 intensitet 3
17038 intensiv 5
17039 intensiva 5
17040 intensivare 1
17041 intensivt 14
17042 intentioner 4
17043 intentionerna 1
17044 inter-etniska 3
17045 interaktiv 3
17046 interaktivitet 2
17047 interaktivitetsnivå 1
17048 interetniska 1
17049 interim 1
17050 interimsavtalen 1
17051 interimsavtalet 4
17052 interimsbetalningar 2
17053 interimsparlament 1
17054 interimspresident 1
17055 interimsråd 2
17056 interimstrukturer 1
17057 interimsåtgärder 1
17058 interinstitutionell 3
17059 interinstitutionella 9
17060 interinstitutionellt 6
17061 intern 14
17062 interna 30
17063 international-socialistiskt 1
17064 internationalisering 1
17065 internationaliseringen 1
17066 internationalistiska 2
17067 internationell 59
17068 internationella 147
17069 internationellt 31
17070 internering 1
17071 interneringar 1
17072 interneringscentra 1
17073 interneringslägret 1
17074 internt 10
17075 interparlamentariska 1
17076 interregionala 4
17077 interregionalt 3
17078 intervenera 2
17079 intervenerar 1
17080 intervention 8
17081 interventioner 5
17082 interventionism 2
17083 interventionskapaciteten 1
17084 interventionsrätt 1
17085 interventionsstödet 1
17086 intervju 2
17087 intervjuades 1
17088 intet 8
17089 intetsägande 1
17090 intill 7
17091 intilliggande 2
17092 intima 1
17093 intimt 4
17094 intog 5
17095 intogs 2
17096 intolerans 5
17097 intoleransen 2
17098 intoleransens 2
17099 intolerant 1
17100 intoleranta 2
17101 intranät 2
17102 intressant 35
17103 intressanta 17
17104 intresse 83
17105 intresseföreningar 1
17106 intresseföreningarna 1
17107 intressekonflikter 2
17108 intressemotsättningar 1
17109 intressen 111
17110 intressena 14
17111 intressenter 1
17112 intressera 4
17113 intresserad 12
17114 intresserade 16
17115 intresserar 10
17116 intresserat 2
17117 intresseregister 1
17118 intresseregistret 2
17119 intressesfärer 1
17120 intresset 10
17121 intrigera 1
17122 intrigerade 1
17123 introducera 1
17124 introducerades 1
17125 introducerat 1
17126 introducerats 2
17127 introduktionskursen 1
17128 introduktionskurser 2
17129 introduktionskurserna 1
17130 intryck 21
17131 intrycket 22
17132 inträdde 1
17133 inträde 5
17134 inträdesbiljett 1
17135 inträffa 17
17136 inträffad 1
17137 inträffade 14
17138 inträffar 15
17139 inträffat 18
17140 intränglingar 1
17141 inträngning 1
17142 inträtt 1
17143 intrång 3
17144 intyg 1
17145 intyga 3
17146 intäkter 11
17147 intäkterna 2
17148 intäktsanalys 1
17149 intäktsbaserade 1
17150 intäktsförluster 1
17151 intåg 1
17152 inuti 2
17153 invaggade 1
17154 invald 1
17155 invandrad 1
17156 invandrade 7
17157 invandrarbefolkningen 1
17158 invandrare 25
17159 invandrares 1
17160 invandrarförläggningar 1
17161 invandrargrupperna 1
17162 invandrarna 6
17163 invandrarnas 2
17164 invandrarpolitik 1
17165 invandring 16
17166 invandringen 7
17167 invandrings- 1
17168 invandringsfientlig 1
17169 invandringsfrågan 1
17170 invandringsfrågorna 1
17171 invandringspolitik 7
17172 invandringspolitiken 2
17173 invandringspolitikens 1
17174 invandringstryck 1
17175 invasion 1
17176 invecklad 2
17177 invecklade 4
17178 invecklar 1
17179 invecklat 2
17180 inventarium 1
17181 inventering 1
17182 inverka 2
17183 inverkan 16
17184 inverkar 5
17185 investera 15
17186 investerade 2
17187 investerar 5
17188 investerare 9
17189 investeraren 1
17190 investerarens 1
17191 investerarna 8
17192 investerarnas 2
17193 investerarskydd 1
17194 investeras 2
17195 investerat 1
17196 investerats 1
17197 investering 7
17198 investeringar 65
17199 investeringarna 14
17200 investeringen 3
17201 investeringsbanken 1
17202 investeringsfonden 1
17203 investeringsfonder 2
17204 investeringsfonderna 1
17205 investeringsfondernas 1
17206 investeringsformer 1
17207 investeringsförmågan 1
17208 investeringskapital 1
17209 investeringskostnader 1
17210 investeringskostnaderna 1
17211 investeringsmöjligheterna 2
17212 investeringsnivån 1
17213 investeringsorgan 1
17214 investeringspolitik 1
17215 investeringspolitiken 1
17216 investeringsslag 1
17217 investeringsspektrumet 1
17218 investeringssyfte 1
17219 investeringsteknikernas 1
17220 investeringstjänstedirektivet 1
17221 investeringstjänster 3
17222 investeringsutgifterna 1
17223 investeringsändamål 2
17224 invid 1
17225 inviga 2
17226 invigd 1
17227 invigdes 2
17228 invigning 2
17229 invigningen 2
17230 invigningsceremonin 1
17231 invigningsfesten 1
17232 invirad 1
17233 invit 1
17234 inviterade 2
17235 involvera 2
17236 involverad 1
17237 involverade 10
17238 involverar 1
17239 involveras 3
17240 invända 2
17241 invändning 5
17242 invändningar 17
17243 invändningen 2
17244 invänta 3
17245 inväntar 1
17246 invånare 21
17247 invånarna 13
17248 invånarnas 1
17249 inälvor 1
17250 inåt 4
17251 inövade 1
17252 iordningställande 1
17253 irakisk 1
17254 irakiska 5
17255 iranske 1
17256 irländarna 1
17257 irländsk 7
17258 irländska 17
17259 irländskt 3
17260 ironi 2
17261 ironisera 1
17262 ironisk 1
17263 ironiska 1
17264 ironiskt 2
17265 irra 1
17266 irrationella 1
17267 irrationellt 1
17268 irreparabla 2
17269 irrgångar 1
17270 irritation 1
17271 irritationsmoment 1
17272 irriterad 4
17273 irriterades 1
17274 irriterar 1
17275 irriterat 1
17276 is 4
17277 iscensatt 1
17278 iscensatte 1
17279 isiga 1
17280 iskalla 1
17281 iskallt 1
17282 isolationism 1
17283 isolera 10
17284 isolerad 1
17285 isolerade 6
17286 isoleras 1
17287 isolerat 4
17288 isolering 7
17289 isoleringseffekter 1
17290 israeler 6
17291 israelerna 6
17292 israelisk 2
17293 israelisk-palestinska 1
17294 israeliska 30
17295 israeliske 1
17296 israeliskt 2
17297 issued 3
17298 istapparna 1
17299 istället 5
17300 isvindar 1
17301 isär 7
17302 it 1
17303 italienarna 2
17304 italiensk 4
17305 italienska 33
17306 italienske 2
17307 italienskt 3
17308 iterationer 1
17309 itu 70
17310 iudice 1
17311 iver 3
17312 ivrig 3
17313 ivriga 1
17314 ivrigt 1
17315 iväg 13
17316 iögonenfallande 2
17317 ja 47
17318 jackärmen 1
17319 jag 3396
17320 jagar 3
17321 jakt 8
17322 jakten 3
17323 jaktområdet 1
17324 jakträtt 1
17325 jamaicanska 1
17326 janela 1
17327 januari 59
17328 januarisessionen 1
17329 janushuvud 1
17330 japaner 1
17331 japanska 1
17332 japanskt 1
17333 jargong 2
17334 jargongen 2
17335 jaså 2
17336 jettons 1
17337 jiddisch 5
17338 jobb 34
17339 jobb-med-framtidsutsikter 1
17340 jobba 4
17341 jobbar 3
17342 jobbat 1
17343 jobben 2
17344 jobbet 4
17345 jobbig 1
17346 joint 1
17347 jojo 1
17348 jojoar 1
17349 jojon 3
17350 jokertecken 5
17351 jokertecknen 2
17352 jokertecknet 1
17353 joniserande 1
17354 jord 14
17355 jordaniska 1
17356 jordbruk 33
17357 jordbrukare 16
17358 jordbrukaren 2
17359 jordbrukares 1
17360 jordbrukarfientliga 1
17361 jordbrukarna 7
17362 jordbrukarnas 3
17363 jordbrukarorganisationer 1
17364 jordbruken 3
17365 jordbruket 36
17366 jordbrukets 7
17367 jordbruks 1
17368 jordbruks- 3
17369 jordbruksaktiviteterna 1
17370 jordbruksavsnittet 1
17371 jordbruksbakgrund 1
17372 jordbruksbefolkningen 1
17373 jordbruksekonomin 1
17374 jordbruksfonden 1
17375 jordbruksfrågornas 1
17376 jordbruksinkomsterna 2
17377 jordbrukskooperativa 1
17378 jordbrukslobbyn 1
17379 jordbruksmarken 1
17380 jordbruksministern 1
17381 jordbruksmodellen 1
17382 jordbruksnäring 1
17383 jordbruksnäringen 2
17384 jordbruksområden 1
17385 jordbruksområdena 2
17386 jordbruksområdenas 1
17387 jordbruksområdet 2
17388 jordbrukspolitik 9
17389 jordbrukspolitiken 25
17390 jordbrukspraxis 1
17391 jordbrukspriserna 1
17392 jordbruksprodukt 1
17393 jordbruksprodukter 4
17394 jordbruksproduktionen 2
17395 jordbruksreformer 1
17396 jordbruksregionerna 1
17397 jordbrukssektorer 1
17398 jordbrukssektorn 12
17399 jordbrukssektorns 1
17400 jordbrukssynpunkt 1
17401 jordbruksutgifterna 1
17402 jordbruksutskott 1
17403 jordbruksutskottet 1
17404 jordbruksutställningar 1
17405 jordbruksverksamhet 1
17406 jordbävningar 1
17407 jordbävningarna 3
17408 jordbävningen 1
17409 jordbävningsdrabbade 1
17410 jordbävningsdramat 1
17411 jordbävningsfara 2
17412 jordbävningssäkra 1
17413 jordbävningsutsatta 1
17414 jorden 10
17415 jordens 8
17416 jordetunnan 1
17417 jordgubbar 1
17418 jordgubbs- 1
17419 jordklotet 1
17420 jordklotets 1
17421 jordluktande 1
17422 jordmån 1
17423 jordnötsformad 1
17424 jordnötssmörglassar 1
17425 jordskalv 1
17426 jordägare 1
17427 journalismen 1
17428 journalist 2
17429 journalisten 10
17430 journalister 8
17431 journalisterna 5
17432 journalisters 1
17433 journalistiska 1
17434 journalists 2
17435 ju 229
17436 jubel 2
17437 jubileumsåret 1
17438 jubla 1
17439 jublande 1
17440 judar 7
17441 judarna 4
17442 judarnas 1
17443 judars 2
17444 jude 6
17445 judegrabbens 1
17446 judeutrotning 1
17447 judisk 3
17448 judiska 6
17449 jugoslaviska 19
17450 jul 2
17451 julen 3
17452 julferien 1
17453 juli 23
17454 julklappar 1
17455 julklappsstämning 1
17456 jumprar 1
17457 jungfrutal 3
17458 juni 40
17459 jure 2
17460 juridisk 14
17461 juridiska 28
17462 juridiskt 16
17463 juris 7
17464 jurisdiktion 7
17465 jurist 1
17466 jurister 3
17467 juristerna 2
17468 juristlingvisterna 1
17469 just 282
17470 justera 3
17471 justerade 1
17472 justerades 6
17473 justerar 2
17474 justeras 3
17475 justering 1
17476 justeringar 4
17477 justeringsfaktor 1
17478 justice 4
17479 justitie- 1
17480 justitiedepartementet 2
17481 justitieminister 1
17482 justitieministern 1
17483 justitieministerns 1
17484 juveler 1
17485 jäkla 2
17486 jämför 6
17487 jämföra 4
17488 jämförande 1
17489 jämföras 2
17490 jämförbar 1
17491 jämförbara 11
17492 jämförbarhet 1
17493 jämförda 1
17494 jämförelse 13
17495 jämförelsen 1
17496 jämförelser 1
17497 jämförelsevis 1
17498 jämförliga 1
17499 jämförligt 1
17500 jämfört 30
17501 jämka 1
17502 jämlik 2
17503 jämlika 2
17504 jämlikar 1
17505 jämlikhet 15
17506 jämlikheten 6
17507 jämlikhetsperspektiv 1
17508 jämlikt 3
17509 jämmer 1
17510 jämn 6
17511 jämna 3
17512 jämnade 2
17513 jämnan 1
17514 jämnt 2
17515 jämnvikten 1
17516 jämsides 2
17517 jämställande 1
17518 jämställd 3
17519 jämställda 2
17520 jämställde 1
17521 jämställdes 1
17522 jämställdhet 28
17523 jämställdheten 8
17524 jämställdhets- 1
17525 jämställdhetsaspekten 2
17526 jämställdhetsdirektiven 1
17527 jämställdhetsfrågor 10
17528 jämställdhetsfrågorna 1
17529 jämställdhetsperspektiv 2
17530 jämställdhetsperspektivet 1
17531 jämställdhetsplanet 1
17532 jämställdhetstänkande 2
17533 jämställdhetstänkandet 1
17534 jämställdhetsutbildning 2
17535 jämställt 1
17536 jämt 4
17537 jämte 2
17538 jämvikt 10
17539 jämvikten 3
17540 järn- 2
17541 järnindustrin 1
17542 järnkrage 1
17543 järnring 1
17544 järnrör 1
17545 järnväg 14
17546 järnvägar 2
17547 järnvägarna 2
17548 järnvägen 6
17549 järnvägens 1
17550 järnvägsföretag 1
17551 järnvägsföretagen 1
17552 järnvägslinjerna 1
17553 järnvägsnät 2
17554 järnvägsnäten 1
17555 järnvägsområde 1
17556 järnvägssektorn 1
17557 järnvägsspår 1
17558 järnvägsövergången 1
17559 järtecken 1
17560 jätte 1
17561 jätteglad 1
17562 jättehårt 1
17563 jättelik 1
17564 jättelikt 1
17565 jätteorder 1
17566 jättestadens 1
17567 jättestor 1
17568 jättestora 2
17569 jättestort 1
17570 jättetankerna 1
17571 jävla 1
17572 k 1
17573 kabarébetonat 1
17574 kabinen 1
17575 kabinett 2
17576 kabinettet 1
17577 kablar 1
17578 kadaver 1
17579 kadmium 4
17580 kadrer 1
17581 kaffe 3
17582 kaffet 2
17583 kafé 2
17584 kajen 1
17585 kaka 1
17586 kakao 1
17587 kakao- 1
17588 kakaoodlarnas 1
17589 kal 1
17590 kala 1
17591 kalender 1
17592 kalkrester 1
17593 kalkylblad 2
17594 kalkylbladsliknande 1
17595 kalkyleras 1
17596 kall 2
17597 kalla 43
17598 kallad 12
17599 kallade 46
17600 kallades 5
17601 kallar 17
17602 kallare 1
17603 kallas 15
17604 kallat 12
17605 kallblodiga 1
17606 kallelse 1
17607 kallelsen 1
17608 kallsvettig 1
17609 kallt 3
17610 kallvattenarter 1
17611 kam 2
17612 kambodjanska 1
17613 kamera 1
17614 kamma 1
17615 kammar 1
17616 kammare 77
17617 kammaren 90
17618 kammarens 9
17619 kammares 4
17620 kamp 28
17621 kampanj 6
17622 kampanjen 3
17623 kampanjer 2
17624 kampen 43
17625 kamrat 2
17626 kamrater 1
17627 kan 2350
17628 kanadensare 1
17629 kanadensisk 1
17630 kanadensiska 3
17631 kanadensiskt 1
17632 kanal 9
17633 kanalen 2
17634 kanaler 6
17635 kanalerna 1
17636 kanderade 1
17637 kandidat 1
17638 kandidater 5
17639 kandidaterna 3
17640 kandidatland 6
17641 kandidatlandstatus 1
17642 kandidatlista 1
17643 kandidatländer 14
17644 kandidatländerna 25
17645 kandidatländernas 8
17646 kandidatprojekten 1
17647 kandidatur 1
17648 kandiderar 2
17649 kanhända 3
17650 kaninen 1
17651 kaniner 1
17652 kaninunge 1
17653 kanoner 2
17654 kanske 200
17655 kansler 2
17656 kanslern 3
17657 kansli 2
17658 kanslichefer 1
17659 kanslierna 1
17660 kanslisekreteraren 1
17661 kant 2
17662 kanten 2
17663 kanter 1
17664 kantonernas 1
17665 kantstött 1
17666 kaos 6
17667 kaotisk 1
17668 kapabel 2
17669 kapacitet 25
17670 kapaciteten 4
17671 kapacitetsbyggnad 1
17672 kapacitetsstöd 1
17673 kapacitetsutveckling 1
17674 kapade 1
17675 kapar 1
17676 kapital 16
17677 kapitalbeskattningen 1
17678 kapitalbildning 1
17679 kapitalet 11
17680 kapitalinkomster 4
17681 kapitalinvesteringstillväxt 1
17682 kapitaliseringsförmåga 1
17683 kapitalistiska 4
17684 kapitalkrav 2
17685 kapitalmarknader 1
17686 kapitalmarknaderna 5
17687 kapitalplaceringar 1
17688 kapitalrörelser 1
17689 kapitalskatt 3
17690 kapitalskatter 1
17691 kapitaltillskott 1
17692 kapitalutnyttjande 1
17693 kapitel 19
17694 kapitelrubrikerna 1
17695 kapitlet 2
17696 kapitulera 1
17697 kapitulerar 1
17698 kapp 2
17699 kapplöpningshaj 1
17700 kapsyler 1
17701 kapten 3
17702 kaptenen 2
17703 kaptener 1
17704 karaff 1
17705 karakteriserade 1
17706 karakteriserar 1
17707 karakteriseringar 1
17708 karakteristisk 1
17709 karakteristiska 1
17710 karakteristiskt 3
17711 karaktär 31
17712 karaktären 8
17713 karaktärer 1
17714 karaktäristisk 1
17715 kareernas 1
17716 karga 2
17717 karikatyr 1
17718 karl 3
17719 karlar 1
17720 karmosinröd 1
17721 karriärer 1
17722 karriärmöjligheter 1
17723 karriärplanering 1
17724 karriärstegen 1
17725 karta 1
17726 kartan 5
17727 kartell- 3
17728 kartellbestämmelserna 1
17729 kartellbildningar 1
17730 karteller 1
17731 kartellförbudet 2
17732 kartellmyndighet 1
17733 kartellrätten 4
17734 kartlägger 1
17735 kartläggning 3
17736 kartonger 1
17737 kartor 2
17738 kasino 2
17739 kaskad 1
17740 kassa 1
17741 kassaapparaten 1
17742 kasserade 3
17743 kassettband 1
17744 kasta 4
17745 kastade 9
17746 kastades 3
17747 kastar 3
17748 kastas 4
17749 kastats 1
17750 kastvapen 1
17751 katalog 4
17752 katalogens 1
17753 katalysator 3
17754 katalytisk 1
17755 katastrof 43
17756 katastrofala 8
17757 katastrofberedskap 1
17758 katastrofdrabbade 3
17759 katastrofen 29
17760 katastrofens 2
17761 katastrofer 34
17762 katastroferna 5
17763 katastrofhjälp 2
17764 katastrofplatsen 1
17765 katastrofprogram 1
17766 katastrofsituation 1
17767 katastrofsituationen 1
17768 katastrofstrategi 1
17769 katastrofstöd 2
17770 kategori 4
17771 kategorier 7
17772 kategorierna 4
17773 kategorifält 3
17774 kategorifältområde 1
17775 kategoriska 1
17776 kategoriskt 1
17777 katolicismen 1
17778 katolik 2
17779 katoliker 3
17780 katolikernas 1
17781 katolska 4
17782 katter 1
17783 kattun 1
17784 kattuntryck 1
17785 kavaj 1
17786 kavaljerer 1
17787 kedja 5
17788 kedjan 5
17789 kedjefångarna 1
17790 kedjorna 1
17791 kejsardömets 1
17792 keltiska 2
17793 kemiindustrins 1
17794 kemikalier 9
17795 kemikaliestrategin 1
17796 kemisk 2
17797 kemiska 13
17798 kg 2
17799 khakishorts 1
17800 khmererna 2
17801 khmerernas 2
17802 kibbutzen 2
17803 kibbutzsjöman 1
17804 kidnappningar 1
17805 kika 1
17806 kil 1
17807 kila 1
17808 kilar 1
17809 kilo 5
17810 kilometer 7
17811 kilowattimme 1
17812 kinderna 1
17813 kindknotor 1
17814 kineser 1
17815 kineserna 3
17816 kinesisk 1
17817 kinesiska 18
17818 kinesiskt 1
17819 kinkig 1
17820 kirurgiskt 1
17821 kisade 1
17822 kittel 1
17823 kitteln 1
17824 kjolarna 1
17825 kl 1
17826 kl. 91
17827 kl.12.00 1
17828 klackar 1
17829 klaga 1
17830 klagade 1
17831 klagan 1
17832 klagar 2
17833 klagat 1
17834 klagoandar 1
17835 klagomål 15
17836 klagomålet 2
17837 klagomålsförfarande 1
17838 klagoskrivelse 1
17839 klagosånger 1
17840 klamrande 1
17841 klandervärt 1
17842 klandras 2
17843 klanen 1
17844 klappa 1
17845 klappjakt 1
17846 klar 42
17847 klara 52
17848 klarade 4
17849 klarades 1
17850 klarar 17
17851 klarare 2
17852 klaras 1
17853 klarast 1
17854 klarat 2
17855 klarats 1
17856 klargjordes 1
17857 klargjort 8
17858 klargör 10
17859 klargöra 25
17860 klargörande 7
17861 klargöranden 3
17862 klargörandet 1
17863 klargöras 4
17864 klargörs 7
17865 klarhet 14
17866 klarheten 1
17867 klarhetens 1
17868 klarlagd 1
17869 klarlagt 1
17870 klarlagts 1
17871 klarlägga 3
17872 klarläggande 4
17873 klarlägganden 2
17874 klarläggandena 1
17875 klarläggandet 1
17876 klarläggas 1
17877 klarsynthet 1
17878 klart 168
17879 klartecken 5
17880 klartext 7
17881 klass 5
17882 klassa 1
17883 klassas 1
17884 klassats 1
17885 klassen 2
17886 klassens 1
17887 klasser 1
17888 klassernas 1
17889 klassificera 3
17890 klassificerar 1
17891 klassificerat 2
17892 klassificering 1
17893 klassificeringen 1
17894 klassificeringsbolagen 1
17895 klassificeringsregister 1
17896 klassificeringssällskapen 4
17897 klassificeringssällskapet 1
17898 klassisk 1
17899 klassiska 4
17900 klassiskt 3
17901 klausul 4
17902 klausulen 2
17903 klausuler 4
17904 klaveret 1
17905 klen 1
17906 klent 1
17907 klev 6
17908 kliande 1
17909 klibbiga 2
17910 klick 2
17911 klient 1
17912 klienter 2
17913 klientilism 1
17914 klimat 12
17915 klimatet 11
17916 klimatfrågor 1
17917 klimatförändring 2
17918 klimatförändringar 5
17919 klimatförändringarna 3
17920 klimatförändringen 2
17921 klimatiska 2
17922 klimatmässiga 1
17923 klimatmönster 1
17924 klimatologiska 2
17925 klimatprotokoll 1
17926 klimatskillnader 1
17927 klingande 1
17928 kliniska 1
17929 kliniskt 1
17930 klippblock 2
17931 klippbranten 1
17932 klippkaos 1
17933 klippstup 1
17934 klippte 1
17935 klirr 1
17936 klirret 1
17937 klistra 1
17938 klistrat 1
17939 kliv 2
17940 kliver 1
17941 kloaklukt 1
17942 klocka 1
17943 klockan 15
17944 klok 6
17945 kloka 2
17946 klokare 2
17947 klokast 1
17948 klokhet 1
17949 klokt 20
17950 klon 1
17951 klorna 1
17952 klotter 1
17953 klumparna 1
17954 klungor 2
17955 klunkar 1
17956 kluven 1
17957 kluvenhet 1
17958 klyfta 2
17959 klyftan 7
17960 klyftor 2
17961 klyftorna 3
17962 klyva 1
17963 klä 2
17964 kläckts 1
17965 klädborste 1
17966 klädd 5
17967 klädda 1
17968 klädde 1
17969 kläder 13
17970 kläderna 2
17971 klädnad 1
17972 klädnader 2
17973 klämde 3
17974 klänning 3
17975 klätt 1
17976 klättra 2
17977 klättrade 2
17978 km 5
17979 knacka 1
17980 knackat 1
17981 knall 1
17982 knallrött 1
17983 knapp 5
17984 knappa 5
17985 knappar 1
17986 knappast 30
17987 knappen 1
17988 knappnålshuvuden 1
17989 knappt 16
17990 knarrar 1
17991 knaster 1
17992 knastrade 1
17993 knep 2
17994 knepiga 1
17995 knipa 1
17996 kniv 2
17997 knivar 2
17998 knivarnas 1
17999 knivhuggen 1
18000 knogande 1
18001 knollrigt 1
18002 knorvig 1
18003 know-how 3
18004 knubbig 1
18005 knuff 1
18006 knussla 1
18007 knuten 6
18008 knutet 3
18009 knutna 9
18010 knutpunkt 1
18011 knutpunkterna 1
18012 knyckte 1
18013 knyta 10
18014 knytas 2
18015 knyter 2
18016 knyts 1
18017 knä 1
18018 knäcka 1
18019 knäckas 1
18020 knäckt 1
18021 knäckte 1
18022 knäna 4
18023 knät 1
18024 knåpat 1
18025 knölar 1
18026 knöt 1
18027 ko 2
18028 ko-affären 1
18029 ko-krisen 1
18030 koalition 3
18031 koalitionen 3
18032 koalitionens 2
18033 koalitionsavtalen 1
18034 koalitionsförhandlingarna 2
18035 koalitionsregering 4
18036 koalitionssamtal 1
18037 kock 1
18038 kockmössa 1
18039 kod 2
18040 koden 3
18041 koder 1
18042 kodifiera 1
18043 kodifierad 3
18044 kodifieras 1
18045 kodifikationen 1
18046 koffertar 1
18047 kofferten 4
18048 koherens 1
18049 koherensen 1
18050 kokade 1
18051 kokhett 1
18052 kokong 1
18053 kokor 1
18054 kokosnötterna 1
18055 kol 1
18056 kol- 1
18057 koldioxid 5
18058 koldioxiden 1
18059 koldioxidutsläppen 1
18060 koleldad 1
18061 kolera 1
18062 kolförrådet 1
18063 kolhög 1
18064 kolja 2
18065 kollaps 1
18066 kollapsa 2
18067 kollega 122
18068 kollegan 26
18069 kollegans 1
18070 kollegas 3
18071 kolleger 266
18072 kollegerna 21
18073 kollegernas 4
18074 kollegers 8
18075 kollegiala 1
18076 kollegialiteten 1
18077 kollegiet 1
18078 kollegium 2
18079 kollegor 32
18080 kollegorna 1
18081 kollegors 4
18082 kollektiv 3
18083 kollektiva 17
18084 kollektivavtal 7
18085 kollektivet 1
18086 kollektivt 2
18087 kollektivtrafik 1
18088 kollektivtrafiken 1
18089 kollisioner 1
18090 kollisionskurs 2
18091 koloni 1
18092 koloniala 2
18093 kolonialdepartementet 1
18094 kolonialdepartementets 1
18095 kolonialism 1
18096 kolonialisterna 1
18097 kolonialmakterna 1
18098 kolonialtiden 1
18099 kolonialtjänsteman 2
18100 kolonialtjänstemännen 1
18101 kolonialtyp 1
18102 kolonier 2
18103 kolonisatörer 3
18104 kolonist 1
18105 kolonisterna 1
18106 koloss 1
18107 kolossala 2
18108 kolossalt 4
18109 kolumn- 2
18110 kolumner 1
18111 kolumnerna 1
18112 kolumnfält 1
18113 kolumnnamn 2
18114 kolumnområden 1
18115 kolumnområdet 1
18116 kolväten 1
18117 kom 141
18118 kombination 7
18119 kombinationen 1
18120 kombinationer 1
18121 kombinera 3
18122 kombinerade 1
18123 kombinerar 3
18124 kombineras 3
18125 kombinerat 1
18126 komedi 1
18127 kometen 1
18128 kometerna 1
18129 komisk 1
18130 komissionen 2
18131 komma 272
18132 kommande 122
18133 kommandon 1
18134 kommandostyrkor 2
18135 kommandot 6
18136 kommas 1
18137 kommen 1
18138 kommendera 1
18139 kommentar 14
18140 kommentarer 36
18141 kommentarerna 4
18142 kommentarsblock 1
18143 kommentatorers 1
18144 kommentera 22
18145 kommenterades 1
18146 kommenterat 1
18147 kommer 1924
18148 kommers 1
18149 kommersiell 5
18150 kommersiella 14
18151 kommersiellt 4
18152 kommission 48
18153 kommissionen 1435
18154 kommissionens 461
18155 kommissionsakt 1
18156 kommissionsdirektoratet 1
18157 kommissionsförslag 1
18158 kommissionskollegiet 1
18159 kommissionsledamot 6
18160 kommissionsledamoten 8
18161 kommissionsledamöter 4
18162 kommissionsledamöterna 3
18163 kommissionsledamöters 1
18164 kommissionsnivå 1
18165 kommissionsordförande 34
18166 kommissionsordföranden 1
18167 kommissionssystemet 1
18168 kommissionstjänsten 1
18169 kommissionär 457
18170 kommissionären 120
18171 kommissionärens 9
18172 kommissionärer 28
18173 kommissionärerna 13
18174 kommissionärernas 2
18175 kommissionärs 1
18176 kommissionärskolleger 1
18177 kommit 92
18178 kommitté 12
18179 kommittédjungel 1
18180 kommittéer 7
18181 kommittéerna 8
18182 kommittéförfarande 2
18183 kommittéförfaranden 6
18184 kommittéförfarandena 2
18185 kommittéförfarandesystemet 2
18186 kommittéförfarandet 16
18187 kommittén 15
18188 kommitténs 1
18189 kommittésystemet 2
18190 kommun 2
18191 kommunal 3
18192 kommunala 7
18193 kommunalparlament 1
18194 kommuner 7
18195 kommunerna 4
18196 kommunfullmäktige 3
18197 kommunicera 1
18198 kommunicerande 1
18199 kommunicerar 1
18200 kommunicerat 1
18201 kommunikation 9
18202 kommunikationen 4
18203 kommunikationer 6
18204 kommunikationerna 1
18205 kommunikations- 1
18206 kommunikationskampanj 1
18207 kommunikationskanaler 2
18208 kommunikationsklyftan 1
18209 kommunikationsmedlen 2
18210 kommunikationsområdet 1
18211 kommunikationsproblemet 1
18212 kommunikationsstrategi 1
18213 kommunikationsteknik 1
18214 kommunikationstekniken 1
18215 kommunikationstjänster 1
18216 kommuniké 1
18217 kommunikéer 1
18218 kommunism 2
18219 kommunismen 1
18220 kommunismens 2
18221 kommunisterna 1
18222 kommunistiska 4
18223 kommunistiskt 2
18224 kommunistpartis 1
18225 kommunistregimerna 1
18226 kommunvalen 1
18227 kompakta 1
18228 kompaniets 1
18229 kompass 1
18230 kompatibelt 2
18231 kompatibla 2
18232 kompensation 17
18233 kompensationer 1
18234 kompensationsfonderna 1
18235 kompensationsåtgärden 1
18236 kompensationsåtgärder 2
18237 kompensationsåtgärderna 2
18238 kompensera 7
18239 kompenserade 1
18240 kompenserades 1
18241 kompenserande 1
18242 kompenserar 3
18243 kompenseras 3
18244 kompenserats 1
18245 kompetens 24
18246 kompetensen 3
18247 kompetenskrav 1
18248 kompetensområden 2
18249 kompetent 8
18250 kompetenta 3
18251 komplement 15
18252 komplementaritet 2
18253 komplementaritetsprinciperna 1
18254 komplett 5
18255 komplettera 23
18256 kompletterad 1
18257 kompletterande 18
18258 kompletterar 5
18259 kompletteras 4
18260 kompletterat 1
18261 komplettering 5
18262 komplex 1
18263 komplexa 5
18264 komplexitet 3
18265 komplexiteten 1
18266 komplext 5
18267 komplicerad 15
18268 komplicerade 11
18269 komplicerat 18
18270 komplikationer 2
18271 komplimang 1
18272 komplimanger 10
18273 komplimentera 1
18274 komplotter 1
18275 komponent 2
18276 komponenten 1
18277 komponenter 8
18278 komponenterna 15
18279 komposteringen 1
18280 kompromettera 1
18281 kompromiss 24
18282 kompromissa 5
18283 kompromissa.§ 1
18284 kompromissarbete 1
18285 kompromissen 5
18286 kompromisser 6
18287 kompromissförslag 4
18288 kompromisslös 1
18289 kompromisslöshet 1
18290 kompromisslösheten 2
18291 kompromisslösning 5
18292 kompromissresolution 1
18293 kompromissresolutionen 4
18294 kompromissrundan 1
18295 kompromisstexten 1
18296 koncentration 14
18297 koncentrationen 6
18298 koncentrationer 7
18299 koncentrationsläger 2
18300 koncentrationslägren 1
18301 koncentrationslägrens 1
18302 koncentrationsprincipen 1
18303 koncentrera 33
18304 koncentrerad 3
18305 koncentrerade 1
18306 koncentrerar 10
18307 koncentreras 7
18308 koncentrerat 5
18309 koncentrerats 1
18310 koncentrisk 1
18311 koncept 10
18312 konceptet 5
18313 koncern 1
18314 koncerner 1
18315 koncis 2
18316 koncisa 1
18317 koncist 2
18318 kondition 1
18319 konfederal 1
18320 konfederation 1
18321 konferens 15
18322 konferensen 21
18323 konferensens 1
18324 konferenserna 3
18325 konfession 1
18326 konfessionslöst 1
18327 konfidentiell 1
18328 konfidentiella 3
18329 konfigurerar 1
18330 konfiskera 1
18331 konfiskerad 1
18332 konfiskerats 1
18333 konflikt 16
18334 konflikten 19
18335 konfliktens 1
18336 konflikter 34
18337 konflikterna 3
18338 konfliktförebyggande 13
18339 konflikthantering 2
18340 konfliktlösning 7
18341 konfliktorsakande 1
18342 konformism 1
18343 konfrontation 1
18344 konfrontationer 1
18345 konfrontationspolitik 1
18346 konfrontera 1
18347 konfronterades 1
18348 konfronteras 7
18349 kongolesisk 1
18350 kongress 1
18351 kongressen 2
18352 kongressmän 1
18353 konjaksglasen 1
18354 konjaksglaset 1
18355 konjunktur 1
18356 konjunkturberoende 1
18357 konjunkturbetingad 1
18358 konjunkturcykeln 1
18359 konjunkturen 3
18360 konjunkturer 1
18361 konjunkturmässiga 1
18362 konjunkturmässigt 1
18363 konjunktursituation 1
18364 konjunktursvängningarna 1
18365 konkret 63
18366 konkreta 104
18367 konkretare 1
18368 konkretaste 1
18369 konkretisera 7
18370 konkretiserar 1
18371 konkretiseras 3
18372 konkretiserats 1
18373 konkretisering 1
18374 konkretiseringar 1
18375 konkurrens 82
18376 konkurrens- 2
18377 konkurrensaspekten 1
18378 konkurrensavgöranden 1
18379 konkurrensbegränsande 2
18380 konkurrensbegränsningar 1
18381 konkurrensbestämmelser 4
18382 konkurrensbestämmelserna 2
18383 konkurrensdebatt 1
18384 konkurrensdebatten 1
18385 konkurrensdomstol 1
18386 konkurrensdugliga 1
18387 konkurrensduglighet 1
18388 konkurrensen 79
18389 konkurrensens 3
18390 konkurrensfriheten 1
18391 konkurrensfrämjande 1
18392 konkurrensfråga 1
18393 konkurrensfrågan 1
18394 konkurrensfrågor 2
18395 konkurrensfrågorna 2
18396 konkurrensfördel 2
18397 konkurrensfördelar 1
18398 konkurrensförfarandet 1
18399 konkurrensförmåga 2
18400 konkurrensförmågan 1
18401 konkurrenshinder 2
18402 konkurrenshämmande 2
18403 konkurrensinitiativen 1
18404 konkurrensinriktad 1
18405 konkurrensjämvikt 1
18406 konkurrenskraft 34
18407 konkurrenskraften 17
18408 konkurrenskraftens 1
18409 konkurrenskraftig 11
18410 konkurrenskraftiga 16
18411 konkurrenskraftigare 2
18412 konkurrenskraftigaste 1
18413 konkurrenskraftigt 2
18414 konkurrenskriterier 1
18415 konkurrenskriterierna 1
18416 konkurrenskultur 3
18417 konkurrenskulturens 1
18418 konkurrenskulturerna 1
18419 konkurrensmedel 1
18420 konkurrensminister 1
18421 konkurrensmyndighet 3
18422 konkurrensmyndigheten 1
18423 konkurrensmyndigheterna 3
18424 konkurrensmyndigheternas 1
18425 konkurrensmyndigheters 1
18426 konkurrensmål 1
18427 konkurrensmöjligheter 1
18428 konkurrensnackdel 1
18429 konkurrensnackdelen 1
18430 konkurrensområdet 3
18431 konkurrensordning 1
18432 konkurrenspakter 1
18433 konkurrenspolitik 20
18434 konkurrenspolitiken 41
18435 konkurrenspolitikens 6
18436 konkurrenspolitisk 1
18437 konkurrenspolitiska 3
18438 konkurrenspolitiskt 2
18439 konkurrensprincipen 3
18440 konkurrenspräglad 1
18441 konkurrensregler 1
18442 konkurrensreglerna 9
18443 konkurrensrelaterade 1
18444 konkurrensrätt 1
18445 konkurrensrätten 6
18446 konkurrensrättens 1
18447 konkurrensrättsliga 1
18448 konkurrenssituationer 1
18449 konkurrensskadlig 1
18450 konkurrensskyddet 2
18451 konkurrensskäl 1
18452 konkurrensstrid 1
18453 konkurrensstörningar 2
18454 konkurrenssvårigheter 1
18455 konkurrenssynpunkt 1
18456 konkurrenstrycket 1
18457 konkurrensutsatt 1
18458 konkurrensutsätta 2
18459 konkurrensutsättning 1
18460 konkurrensutsättningar 1
18461 konkurrensutsättningen 1
18462 konkurrensverken 1
18463 konkurrensvillkor 5
18464 konkurrensvillkoren 7
18465 konkurrensvänligare 1
18466 konkurrensärenden 2
18467 konkurrent 2
18468 konkurrenter 7
18469 konkurrentländer 1
18470 konkurrera 11
18471 konkurrerar 1
18472 konkurs 3
18473 konkurser 5
18474 konkursfond 1
18475 konsekvens 16
18476 konsekvensen 3
18477 konsekvenser 64
18478 konsekvenserna 36
18479 konsekvensutredning 2
18480 konsekvensutredningar 2
18481 konsekvensutredningarnas 1
18482 konsekvent 27
18483 konsekventa 9
18484 konsensus 2
18485 konsert 1
18486 konserten 1
18487 konservativa 13
18488 konservativas 1
18489 konserver 1
18490 konsolidera 1
18491 konsoliderade 1
18492 konsoliderar 1
18493 konsoliderat 1
18494 konsolidering 5
18495 konsolideringen 3
18496 konsolideringsprogram 1
18497 konsortierna 1
18498 konspirationer 1
18499 konst 5
18500 konstant 4
18501 konstatera 69
18502 konstaterade 4
18503 konstaterades 2
18504 konstaterande 4
18505 konstaterandet 2
18506 konstaterar 12
18507 konstateras 4
18508 konstaterat 7
18509 konstaterats 1
18510 konsten 1
18511 konstfullt 1
18512 konstföremål 1
18513 konstgjord 2
18514 konstgjorda 1
18515 konstgjort 1
18516 konstgrepp 1
18517 konstgödsel 1
18518 konstig 1
18519 konstiga 2
18520 konstigt 6
18521 konstituera 1
18522 konstituerades 1
18523 konstitution 5
18524 konstitutionell 4
18525 konstitutionella 23
18526 konstitutionen 1
18527 konstitutivt 1
18528 konstkommittén 1
18529 konstkritikern 1
18530 konstlade 1
18531 konstlat 1
18532 konstlöst 1
18533 konstmuseum 1
18534 konstnären 1
18535 konstnärer 5
18536 konstnärerna 4
18537 konstnärers 4
18538 konstnärliga 3
18539 konstruera 6
18540 konstruerades 1
18541 konstruerat 1
18542 konstruerats 1
18543 konstruktion 9
18544 konstruktionen 1
18545 konstruktioner 1
18546 konstruktionsarbete 1
18547 konstruktionsarbetet 5
18548 konstruktiv 9
18549 konstruktiva 15
18550 konstruktivt 12
18551 konstruktören 1
18552 konstruktörerna 1
18553 konststycken 1
18554 konstverk 1
18555 konsultationer 3
18556 konsultbasis 1
18557 konsulter 1
18558 konsulterande 1
18559 konsulteras 1
18560 konsument 2
18561 konsumenten 16
18562 konsumenten-medborgaren 1
18563 konsumenter 16
18564 konsumenterna 32
18565 konsumenternas 25
18566 konsumenters 1
18567 konsumentfrågor 20
18568 konsumentförtroende 1
18569 konsumentorganisationen 1
18570 konsumentpolitik 4
18571 konsumentpolitisk 1
18572 konsumentrelaterad 1
18573 konsumenträtten 1
18574 konsumentskydd 11
18575 konsumentskyddet 6
18576 konsumentskyddsorganisationerna 1
18577 konsumenttillvänt 1
18578 konsumentvaror 1
18579 konsumentvänligt 1
18580 konsumeras 1
18581 konsumtion 4
18582 konsumtionen 2
18583 kontakt 19
18584 kontaktade 1
18585 kontaktat 3
18586 kontakten 5
18587 kontakter 23
18588 kontakterna 5
18589 kontamination 1
18590 kontaminerade 1
18591 kontanter 1
18592 kontexten 1
18593 kontinent 9
18594 kontinentala 3
18595 kontinentaleuropéerna 1
18596 kontinentalt 1
18597 kontinenten 7
18598 kontinentens 3
18599 kontinenter 1
18600 kontinenterna 1
18601 kontinents 2
18602 kontinuerlig 3
18603 kontinuerligt 4
18604 kontinuitet 3
18605 kontinuiteten 3
18606 kontor 10
18607 kontoren 1
18608 kontoret 2
18609 kontorslokaler 1
18610 kontrahenterna 1
18611 kontrakt 9
18612 kontraktet 2
18613 kontrakts- 1
18614 kontraktsramar 1
18615 kontraktsåtagande 1
18616 kontraproduktiv 1
18617 kontraproduktivt 2
18618 kontrast 3
18619 kontrasten 1
18620 kontraster 1
18621 kontrasterar 1
18622 kontroll 119
18623 kontroll- 2
18624 kontrollanterna 1
18625 kontrollapparat 1
18626 kontrollen 32
18627 kontroller 44
18628 kontrollera 44
18629 kontrollerad 5
18630 kontrollerade 3
18631 kontrollerades 1
18632 kontrollerar 9
18633 kontrolleras 19
18634 kontrollerat 1
18635 kontrollerbara 1
18636 kontrollerna 6
18637 kontrollfunktion 1
18638 kontrollförfarande 1
18639 kontrollförfaranden 2
18640 kontrollförfarandet 1
18641 kontrollmakt 1
18642 kontrollmakten 1
18643 kontrollmedlen 1
18644 kontrollmekanismer 3
18645 kontrollmyndighet 1
18646 kontrollmyndigheterna 1
18647 kontrollmöjlighet 1
18648 kontrollmöjligheter 3
18649 kontrollnormerna 1
18650 kontrollområdet 1
18651 kontrollorgan 2
18652 kontrollprocessen 1
18653 kontrollprogram 1
18654 kontrollprogrammen 1
18655 kontrollrättigheter 1
18656 kontrollstyrka 1
18657 kontrollsystem 2
18658 kontrollsystemet 1
18659 kontrollsystemets 1
18660 kontrolluppdrag 1
18661 kontrollverksamheten 1
18662 kontrolläger 1
18663 kontrollåtgärder 2
18664 kontrovers 2
18665 kontroversen 2
18666 kontroverser 3
18667 kontroversiell 4
18668 kontroversiella 2
18669 kontroversiellt 4
18670 konturlösa 1
18671 konungariket 1
18672 konvenansflagg 1
18673 konvent 2
18674 konventet 3
18675 konvention 23
18676 konventionella 2
18677 konventionen 37
18678 konventionens 2
18679 konventioner 12
18680 konventionerna 1
18681 konventionsinstrumenten 1
18682 konventionsnivå 1
18683 konvergens 20
18684 konvergensen 9
18685 konvergenskriterier 6
18686 konvergenskriterierna 3
18687 konvergenskriterium 2
18688 konvergensperspektiv 1
18689 konvergensprocess 1
18690 konvergensprogrammen 1
18691 konvergensstrategi 1
18692 konvergensstrategier 1
18693 konvergensstrategin 1
18694 konvergering 1
18695 konvergeringsprocess 1
18696 konversation 1
18697 konversationen 1
18698 konverserade 1
18699 konvertera 4
18700 konverterade 2
18701 konverteras 3
18702 kooperationens 1
18703 kooperativ 1
18704 kooperativa 1
18705 kopia 3
18706 kopian 1
18707 kopiera 4
18708 kopierade 3
18709 kopierar 5
18710 kopieras 2
18711 kopiering 4
18712 kopieringsrätten 1
18713 kopieringsskyddet 1
18714 kopior 3
18715 kopp 1
18716 koppar 1
18717 kopparbrunt 1
18718 koppen 1
18719 koppla 4
18720 kopplad 3
18721 kopplas 5
18722 kopplat 2
18723 kopplats 1
18724 koppling 8
18725 kopplingarna 1
18726 kopplingen 4
18727 kor 1
18728 kor. 1
18729 korgar 1
18730 korken 1
18731 korna 1
18732 korporatism 1
18733 korpsvart 1
18734 korpus 1
18735 korrekt 44
18736 korrekta 11
18737 korrektare 2
18738 korrekthet 1
18739 korrespondens 1
18740 korrespondent 1
18741 korrespondenten 1
18742 korrespondenter 1
18743 korridoren 1
18744 korridorer 3
18745 korridorerna 1
18746 korridorernas 1
18747 korrigerande 1
18748 korrigeras 1
18749 korrugerad 1
18750 korrumpera 1
18751 korrumperat 2
18752 korrupt 1
18753 korrupta 1
18754 korruption 14
18755 korruptionen 9
18756 korruptionsaffärer 3
18757 korruptionsdömt 1
18758 korruptionsskandal 1
18759 korruptionsskandalerna 1
18760 kors 2
18761 korsade 2
18762 korsar 1
18763 korseld 1
18764 korselden 1
18765 korset 2
18766 korsett 1
18767 korsfråga 4
18768 korslagda 1
18769 korsriddarna 1
18770 kort 132
18771 korta 17
18772 kortare 6
18773 kortas 3
18774 kortaste 1
18775 korten 2
18776 kortet 7
18777 kortets 3
18778 kortfattad 1
18779 kortfattat 2
18780 korthet 3
18781 kortlek 1
18782 kortlivad 1
18783 kortsiktig 2
18784 kortsiktiga 4
18785 kortsiktighet 2
18786 kortsiktigt 2
18787 kortsnaggade 1
18788 kortvarig 1
18789 kortväxt 2
18790 korvar 1
18791 koscherlunch 2
18792 koschermat 2
18793 koschersmörgåsar 1
18794 kosovanska 1
18795 kosovoalbaner 6
18796 kosovoalbanerna 3
18797 kosovoalbanska 2
18798 kosta 4
18799 kostade 5
18800 kostar 14
18801 kostat 2
18802 kosthållning 1
18803 kostnad 14
18804 kostnaden 26
18805 kostnader 59
18806 kostnaderna 61
18807 kostnads 1
18808 kostnads- 1
18809 kostnads-intäktsanalys 1
18810 kostnads-intäktsanalysen 1
18811 kostnads-nytto-analys 1
18812 kostnadsbefrielse 1
18813 kostnadsbefrielsen 3
18814 kostnadseffektiv 2
18815 kostnadseffektiva 2
18816 kostnadseffektivt 1
18817 kostnadselementet 1
18818 kostnadsfri 3
18819 kostnadsfria 1
18820 kostnadsfritt 1
18821 kostnadsfördelningen 1
18822 kostnadsinflation 1
18823 kostnadsintensiv 1
18824 kostnadsintensivt 1
18825 kostnadskontroll 1
18826 kostnadspolicy 1
18827 kostnadssystem 4
18828 kostnadstäckande 1
18829 kostnadstäckning 1
18830 kostnadsuppskattning 1
18831 kostnadsutvecklingen 1
18832 kostsam 1
18833 kostsamma 1
18834 kostsamt 3
18835 kostym 1
18836 kostymen 1
18837 kovändning 1
18838 krafsar 1
18839 kraft 83
18840 kraften 11
18841 krafter 16
18842 krafterna 4
18843 krafters 1
18844 kraftfull 6
18845 kraftfulla 10
18846 kraftfullare 2
18847 kraftfullt 16
18848 kraftig 15
18849 kraftiga 8
18850 kraftigare 4
18851 kraftigaste 1
18852 kraftigt 31
18853 kraftmätning 1
18854 kraftnät 1
18855 krafttag 3
18856 kraftåtgärder 1
18857 kragar 1
18858 kragen 1
18859 kramade 1
18860 kramat 1
18861 krampen 1
18862 kran 1
18863 kranarna 1
18864 krasande 1
18865 kraschade 1
18866 kraschat 1
18867 krasst 1
18868 krav 119
18869 kravallpoliser 1
18870 kraven 37
18871 kravet 31
18872 kravla 1
18873 kreativ 2
18874 kreativa 4
18875 kreativitet 1
18876 kreativiteten 3
18877 kreativt 1
18878 kreatörer 1
18879 krediter 1
18880 krediterna 1
18881 kreditinstitut 1
18882 kreditvärdighet 2
18883 kreditvärdighetsskala 1
18884 kretensare 1
18885 krets 1
18886 kretsar 3
18887 kretsat 1
18888 kretsen 2
18889 kretslopp 3
18890 krig 46
18891 kriga 2
18892 krigare 1
18893 krigat 1
18894 krigen 2
18895 kriget 30
18896 krigföring 2
18897 krigisk 2
18898 krigsekonomi 1
18899 krigsfartyg 1
18900 krigsflyktingar 1
18901 krigsfångar 1
18902 krigsförbrytardomstolen 1
18903 krigsförbrytare 1
18904 krigsförbrytartribunalen 4
18905 krigsförbrytelser 1
18906 krigsförklaring 1
18907 krigshandlingar 1
18908 krigshandlingarna 1
18909 krigsherrarna 1
18910 krigshärjade 1
18911 krigsivrare 1
18912 krigskonstens 1
18913 krigskorrespondenten 1
18914 krigsmaskin 1
18915 krigsmateriel 1
18916 krigsmålad 1
18917 krigspropagandan 1
18918 krigssituationer 1
18919 krigsskador 1
18920 krigsslutet 1
18921 krigsterminalen 1
18922 krigsutbrott 1
18923 krigsåren 1
18924 kriminalisera 2
18925 kriminaliseras 1
18926 kriminalitet 8
18927 kriminalitetsbekämpning 1
18928 kriminalpolitik 1
18929 kriminalvården 1
18930 kriminell 1
18931 kriminella 5
18932 kriminellt 1
18933 kring 51
18934 kringgå 3
18935 kringgående 2
18936 kringgår 1
18937 kringgås 1
18938 kringirrande 1
18939 kringliggande 1
18940 kringskuren 1
18941 kringskuret 1
18942 kringspridda 1
18943 kringströvanden 1
18944 kringvärvd 1
18945 kringvärvde 1
18946 kris 19
18947 krisbildningarna 1
18948 kriscenter 1
18949 krisen 11
18950 krisens 1
18951 kriser 13
18952 krisförebyggande 1
18953 krisförordning 1
18954 krishantering 9
18955 krishanteringsplanerna 1
18956 krisläge 1
18957 krisläget 1
18958 krismedvetande 2
18959 krismöte 1
18960 krisområde 1
18961 krisområden 1
18962 krisperioden 1
18963 krisregionen 1
18964 krissituationen 1
18965 krissituationer 1
18966 krisstyrningsåtgärderna 1
18967 kristallklara 2
18968 kristdemokrater 20
18969 kristdemokraterna 5
18970 kristdemokraternas 1
18971 kristdemokratisk 1
18972 kristdemokratiska 1
18973 kristdemokratiske 1
18974 kristendom 1
18975 kristendomens 1
18976 kristna 1
18977 kritan 4
18978 kriterier 38
18979 kriterierna 8
18980 kriteriet 1
18981 kriterium 1
18982 kritik 28
18983 kritiken 10
18984 kritiker 2
18985 kritisera 18
18986 kritiserade 1
18987 kritiserades 1
18988 kritiserar 10
18989 kritiseras 3
18990 kritiserat 3
18991 kritiserats 1
18992 kritisk 20
18993 kritiska 17
18994 kritiskt 8
18995 kroater 1
18996 krocka 1
18997 krog 1
18998 krok 1
18999 krokar 2
19000 krokig 1
19001 krom 3
19002 krombrickor 1
19003 kromen 1
19004 kronan 1
19005 kronjuvelen 1
19006 kropp 8
19007 kroppar 1
19008 kroppen 4
19009 kroppens 1
19010 kropps 1
19011 kroppsbyggnad 1
19012 kroppslösa 1
19013 kroppsrytm 1
19014 kroppstemperatur 1
19015 krossa 1
19016 krossar 1
19017 krukpalm 1
19018 krukskärva 1
19019 krumryggad 1
19020 krutdurk 1
19021 krutet 1
19022 krutröken 1
19023 kryddgården 1
19024 kryllar 1
19025 krympande 1
19026 kryphål 4
19027 kryphålen 1
19028 kryssa 1
19029 kryssningen 2
19030 kräftgång 1
19031 kränka 2
19032 kränkande 1
19033 kränker 5
19034 kränkning 9
19035 kränkningar 16
19036 kränkningarna 10
19037 kränks 5
19038 kränkt 1
19039 kränkta 1
19040 kränkts 1
19041 kräva 62
19042 krävande 7
19043 krävas 8
19044 krävde 6
19045 krävdes 7
19046 kräver 130
19047 krävs 147
19048 krävt 10
19049 krävts 2
19050 krångel 1
19051 krångla 1
19052 krånglar 1
19053 krånglig 1
19054 krångliga 1
19055 krökte 1
19056 krönas 1
19057 krönikör 2
19058 kröp 1
19059 kubanerna 1
19060 kubanernas 1
19061 kubansk 1
19062 kubanska 3
19063 kubikmeter 2
19064 kudde 1
19065 kudden 1
19066 kula 2
19067 kuliss 1
19068 kulisserna 4
19069 kullar 1
19070 kulle 1
19071 kullerstensgatan 1
19072 kullkasta 1
19073 kullkastar 1
19074 kullvräkt 1
19075 kulmen 1
19076 kulminerade 1
19077 kulor 1
19078 kultiverad 1
19079 kultur 62
19080 kultur- 2
19081 kulturaktiviteter 1
19082 kulturanslag 1
19083 kulturarbetare 1
19084 kulturarv 7
19085 kulturarvet 2
19086 kulturell 19
19087 kulturella 26
19088 kulturella-historiska 1
19089 kulturellt 15
19090 kulturen 23
19091 kulturens 4
19092 kulturer 4
19093 kulturerna 1
19094 kulturform 1
19095 kulturförändring 1
19096 kulturhistoriskt 1
19097 kulturindustripolitik 1
19098 kulturområde 4
19099 kulturområdet 1
19100 kulturpolitik 5
19101 kulturpolitikens 1
19102 kulturpolitiska 1
19103 kulturprogram 2
19104 kulturprogrammet 1
19105 kulturresurserna 1
19106 kultursektorn 4
19107 kultursektors 1
19108 kulturservice 1
19109 kulturskillnader 1
19110 kulturutskottet 1
19111 kumulativa 3
19112 kumulativt 1
19113 kumuleringen 1
19114 kund 2
19115 kunde 214
19116 kunden 3
19117 kundens 1
19118 kunder 9
19119 kunderna 4
19120 kundernas 3
19121 kundkretsen 1
19122 kundorderformat 1
19123 kundorientering 1
19124 kundrelation 1
19125 kundvagnen 1
19126 kundvänliga 1
19127 kung 1
19128 kungariket 33
19129 kungarikets 12
19130 kungars 1
19131 kungen 1
19132 kungliga 1
19133 kungssportfiskare 1
19134 kunna 624
19135 kunnande 7
19136 kunnat 107
19137 kunnig 1
19138 kunnigt 1
19139 kunskap 26
19140 kunskapen 4
19141 kunskapens 2
19142 kunskaper 10
19143 kunskaperna 3
19144 kunskapsbaserad 3
19145 kunskapsbristen 1
19146 kunskapsdrivna 1
19147 kunskapsekonomi 2
19148 kunskapsekonomin 5
19149 kunskapsmässig 1
19150 kunskapsområdena 1
19151 kunskapssamhälle 4
19152 kunskapssamhället 7
19153 kunskapsspridning 1
19154 kunskapsträning 1
19155 kunskapsuppbyggnad 1
19156 kunskapsutveckling 1
19157 kunskapsöverföring 1
19158 kurade 1
19159 kurder 1
19160 kurdiska 1
19161 kurs 4
19162 kursen 2
19163 kurser 1
19164 kurserna 1
19165 kursriktning 1
19166 kursändring 3
19167 kurva 2
19168 kusinen 1
19169 kusiner 1
19170 kusligt 1
19171 kust 7
19172 kust- 1
19173 kustbefolkningarnas 1
19174 kustbevakningen 1
19175 kustbevakningskårer 1
19176 kustbevakningsstyrka 1
19177 kusten 19
19178 kustens 1
19179 kuster 6
19180 kusterna 8
19181 kusternas 1
19182 kustfiskebåtar 1
19183 kustfisket 1
19184 kusthamnarna 1
19185 kustland 1
19186 kustlinje 2
19187 kustmyndigheter 2
19188 kustmyndigheternas 1
19189 kustneger 1
19190 kustnära 2
19191 kustområden 9
19192 kustområdena 3
19193 kustregioner 1
19194 kustregionerna 2
19195 kuststad 1
19196 kustvakter 1
19197 kustvatten 2
19198 kustvattnen 1
19199 kuvert 1
19200 kval 1
19201 kvalificera 2
19202 kvalificerad 20
19203 kvalificerade 8
19204 kvalificerat 3
19205 kvalifikationer 3
19206 kvalitativ 6
19207 kvalitativa 7
19208 kvalitativt 8
19209 kvalitet 54
19210 kvaliteten 34
19211 kvaliteter 2
19212 kvalitetsbevarande 1
19213 kvalitetsförbättringar 1
19214 kvalitetsförluster 1
19215 kvalitetsförsämring 1
19216 kvalitetsgaranti 1
19217 kvalitetskontroll 1
19218 kvalitetskrav 1
19219 kvalitetskraven 1
19220 kvalitetskriterier 1
19221 kvalitetsmätningen 1
19222 kvalitetsmålen 1
19223 kvalitetsnivå 1
19224 kvalitetsnormer 3
19225 kvalitetsprojekt 1
19226 kvalitetssprång 1
19227 kvalitén 1
19228 kvalmigt 1
19229 kvantifierade 3
19230 kvantifieras 1
19231 kvantifierbara 4
19232 kvantitativ 3
19233 kvantitativa 9
19234 kvantitativt 3
19235 kvantitet 3
19236 kvantiteter 1
19237 kvantitetsgränser 1
19238 kvantitetshantering 1
19239 kvantitetshanteringen 1
19240 kvar 80
19241 kvarhängande 1
19242 kvarhålla 1
19243 kvarhållandena 1
19244 kvarhåller 1
19245 kvarhölls 1
19246 kvarleva 1
19247 kvarnsten 1
19248 kvarstad 1
19249 kvarstå 1
19250 kvarstår 10
19251 kvarstått 1
19252 kvartalet 1
19253 kvarter 8
19254 kvarteren 1
19255 kvarvarande 3
19256 kvasten 1
19257 kvastkäppen 1
19258 kvav 1
19259 kvavt 1
19260 kvestor 1
19261 kvestorer 3
19262 kvestorerna 9
19263 kvestorernas 1
19264 kvestorskollegiet 1
19265 kvickhet 1
19266 kvicksilver 6
19267 kvickt 1
19268 kvinna 25
19269 kvinnan 8
19270 kvinnans 4
19271 kvinnfolk 1
19272 kvinnlig 6
19273 kvinnliga 20
19274 kvinnlighet 1
19275 kvinnligt 2
19276 kvinnodagen 5
19277 kvinnofrågan 1
19278 kvinnogrupperna 1
19279 kvinnohandel 2
19280 kvinnokonferensen 1
19281 kvinnoprogrammet 2
19282 kvinnor 182
19283 kvinnorepresentationen 1
19284 kvinnorna 46
19285 kvinnornas 23
19286 kvinnors 45
19287 kvinnorörelsens 1
19288 kvinnoutskott 1
19289 kvinnoutskottet 1
19290 kvinnspersoner 1
19291 kvistar 1
19292 kvitt 2
19293 kvitterade 1
19294 kvot 10
19295 kvoten 3
19296 kvoter 17
19297 kvoterad 1
19298 kvotering 8
19299 kvoteringar 1
19300 kvoteringspolitik 1
19301 kvoteringspåföljder 1
19302 kvoterna 2
19303 kvotflyktingar 1
19304 kvotsystemet 1
19305 kväll 40
19306 kvällar 3
19307 kvällarna 2
19308 kvällen 11
19309 kvällens 4
19310 kvällningen 1
19311 kvällsmat 1
19312 kvällsmöte 1
19313 kväva 4
19314 kväve 1
19315 kyckling 4
19316 kycklingar 2
19317 kycklingarna 1
19318 kycklingen 1
19319 kyla 3
19320 kylan 3
19321 kyliga 2
19322 kyligt 1
19323 kylskåpet 2
19324 kylstela 1
19325 kypare 1
19326 kyrkan 1
19327 kyrkans 2
19328 kyrkdörren 1
19329 kyrkogård 1
19330 kyrkorna 3
19331 kyrkpiano 1
19332 kyss 1
19333 kyssa 1
19334 kysste 1
19335 käbbel 1
19336 käbblade 1
19337 käckt 1
19338 käll- 1
19339 källa 15
19340 källan 5
19341 källare 1
19342 källaren 1
19343 källformat 1
19344 källor 7
19345 källorna 2
19346 kämpa 8
19347 kämpade 2
19348 kämpar 7
19349 kämpat 3
19350 känd 7
19351 kända 13
19352 kände 39
19353 kändes 14
19354 känn 2
19355 känna 38
19356 kännas 1
19357 kännbar 1
19358 kännbart 1
19359 kännedom 9
19360 kännedomen 1
19361 känner 164
19362 kännetecken 1
19363 känneteckna 2
19364 kännetecknade 1
19365 kännetecknades 2
19366 kännetecknande 1
19367 kännetecknar 1
19368 kännetecknas 7
19369 kännetecknat 1
19370 känns 3
19371 känsla 22
19372 känslan 12
19373 känslans 1
19374 känslig 23
19375 känsliga 17
19376 känsligare 2
19377 känsligaste 3
19378 känslighet 5
19379 känsligt 7
19380 känslokall 1
19381 känslokalla 1
19382 känsloladdad 1
19383 känslomässiga 2
19384 känslomässigt 1
19385 känslor 10
19386 känslotänkande 1
19387 känt 22
19388 känts 1
19389 käpp 1
19390 käpprakt 1
19391 kär 2
19392 kära 111
19393 käre 2
19394 kärl 1
19395 kärlek 4
19396 kärleken 4
19397 kärna 6
19398 kärnaktivitet 1
19399 kärnan 8
19400 kärnenergisäkerhet 6
19401 kärnenergisäkerhetsfördragen 1
19402 kärnenergiäkerhet 1
19403 kärnfission 1
19404 kärnforskning 1
19405 kärnfrågan 2
19406 kärnfrågor 1
19407 kärnfusion 1
19408 kärnkatastrofer 1
19409 kärnkraft 5
19410 kärnkraften 1
19411 kärnkraftens 1
19412 kärnkraftsanläggningar 3
19413 kärnkraftsanläggningarna 1
19414 kärnkraftsolycka 1
19415 kärnkraftsolyckor 1
19416 kärnkraftsområdet 1
19417 kärnkraftsplanerna 1
19418 kärnkraftsprogram 1
19419 kärnkraftsreaktorer 1
19420 kärnkraftssäkerhet 1
19421 kärnkraftsverk 1
19422 kärnkraftverk 7
19423 kärnkraftverken 1
19424 kärnområden 1
19425 kärnprinciper 1
19426 kärnprinciperna 1
19427 kärnproblemen 1
19428 kärnpunkt 1
19429 kärnpunkten 2
19430 kärnpunkter 1
19431 kärnstrålningskontroller 1
19432 kärnsäkerhet 3
19433 kärnteknik 2
19434 kärnuppgifter 1
19435 kärnuppgifterna 1
19436 kärnvapen 6
19437 kärnvapenspridning 1
19438 kärnvapenteknik 1
19439 kärnvapenutveckling 1
19440 kärnverksamhet 1
19441 kärran 2
19442 kål 3
19443 kålhuven 1
19444 kånkande 1
19445 kår 1
19446 kåren 2
19447 kårer 1
19448 kö 2
19449 köat 1
19450 köer 1
19451 kök 2
19452 köket 11
19453 köksbiträde 2
19454 köksbordet 2
19455 köksstolen 1
19456 köl 3
19457 kölar 1
19458 köld 3
19459 köldbeständigheten 1
19460 köldgränsen 1
19461 kölvattnet 1
19462 kön 12
19463 könen 15
19464 könens 1
19465 könet 1
19466 könsapartheid 1
19467 könsdiskriminering 1
19468 könsfrågor 1
19469 könsfördelning 2
19470 könsförändringar 1
19471 könsgrundade 1
19472 könsidentiteter 1
19473 könskvotering 5
19474 könsorgan 1
19475 könsrelaterad 1
19476 könsrelaterade 1
19477 könsspecifika 1
19478 köp 1
19479 köpa 5
19480 köpare 1
19481 köpas 1
19482 köpenskap 1
19483 köper 4
19484 köpet 4
19485 köpkraft 1
19486 köpkraften 1
19487 köpmans 1
19488 köps 1
19489 köpslagningslogik 1
19490 köpslå 1
19491 köpt 3
19492 köpte 6
19493 kör 8
19494 köra 5
19495 köras 5
19496 körde 5
19497 kördes 1
19498 körförbud 1
19499 körning 1
19500 körningen 1
19501 körningsfel 1
19502 körs 3
19503 körsbärs- 1
19504 kört 4
19505 körtid 1
19506 körtidsfunktioner 1
19507 kött 2
19508 kött- 1
19509 köttkrig 1
19510 köttprodukter 1
19511 köttskiva 1
19512 l 1
19513 l'Etat 2
19514 l'Europe 1
19515 l'eau 1
19516 la 8
19517 laboratorier 1
19518 laboratorium 2
19519 laborerar 2
19520 labourkolleger 1
19521 labourledamöterna 1
19522 labourledamöternas 1
19523 labours 2
19524 labradoren 1
19525 labyrint 1
19526 lackstång 1
19527 lackstången 1
19528 laddat 2
19529 lade 48
19530 lades 15
19531 lag 19
19532 laga 2
19533 lagade 2
19534 lagar 30
19535 lagarna 5
19536 lagbrott 1
19537 lagd 1
19538 lagen 19
19539 lagenligt 1
19540 lagens 2
19541 lager 6
19542 lagerhus 2
19543 lagerkrans 1
19544 laget 6
19545 lagförslag 6
19546 lagförslaget 2
19547 lagkränkning 1
19548 laglig 1
19549 lagliga 6
19550 laglighet 2
19551 lagligheten 1
19552 lagligt 8
19553 lagmängden 1
19554 lagom 1
19555 lagra 3
19556 lagrade 2
19557 lagrar 1
19558 lagras 1
19559 lagret 1
19560 lagring 1
19561 lagringskapacitet 1
19562 lags 1
19563 lagstadgad 1
19564 lagstadgade 2
19565 lagstifta 7
19566 lagstiftande 19
19567 lagstiftar 5
19568 lagstiftare 1
19569 lagstiftarna 2
19570 lagstiftat 2
19571 lagstiftning 124
19572 lagstiftningar 2
19573 lagstiftningen 59
19574 lagstiftningens 1
19575 lagstiftnings- 1
19576 lagstiftningsarbete 1
19577 lagstiftningsarbetet 6
19578 lagstiftningscykel 1
19579 lagstiftningsfrågor 1
19580 lagstiftningsförfarande 2
19581 lagstiftningsförfarandet 4
19582 lagstiftningsförslag 6
19583 lagstiftningsinitiativ 2
19584 lagstiftningsinstrument 1
19585 lagstiftningsmängd 1
19586 lagstiftningsområden 2
19587 lagstiftningsperioden 1
19588 lagstiftningsprocess 1
19589 lagstiftningsprocessen 5
19590 lagstiftningsprogram 9
19591 lagstiftningsprogrammet 8
19592 lagstiftningsramen 1
19593 lagstiftningsreformen 1
19594 lagstiftningsresolutionen 10
19595 lagstiftningsresolutionerna 2
19596 lagstiftningsåtgärder 5
19597 lagt 101
19598 lagtext 2
19599 lagtexten 1
19600 lagtexter 1
19601 lagtexterna 1
19602 lagts 49
19603 lagändringar 1
19604 laissez 1
19605 lamaismen 1
19606 lambala-talande 1
19607 lamm 1
19608 lampa 1
19609 lampor 1
19610 lamporna 1
19611 lamslagen 1
19612 land 266
19613 landades 1
19614 landar 1
19615 landas 2
19616 landat 1
19617 landats 1
19618 landet 72
19619 landets 21
19620 landgränserna 2
19621 landminor 5
19622 landmärke 1
19623 landning 1
19624 landningen 1
19625 landningsbanan 1
19626 landområde 1
19627 landområden 1
19628 landpermission 2
19629 landremsan 1
19630 lands 15
19631 landsatte 3
19632 landsbruket 1
19633 landsbygd 3
19634 landsbygden 67
19635 landsbygdens 28
19636 landsbygdsbefolkningarna 1
19637 landsbygdsbefolkningen 1
19638 landsbygdskommuners 1
19639 landsbygdsområde 1
19640 landsbygdsområden 10
19641 landsbygdsområdena 3
19642 landsbygdsområdet 9
19643 landsbygdsområdets 1
19644 landsbygdspolitiken 1
19645 landsbygdsproblem 1
19646 landsbygdsregion 1
19647 landsbygdsregioner 2
19648 landsbygdsregionerna 2
19649 landsbygdsstrukturens 1
19650 landsbygdsturism 1
19651 landsbygdsutveckling 13
19652 landsbygdsutvecklingen 2
19653 landsbygdsutvecklingens 1
19654 landsflykten 1
19655 landsförvisning 2
19656 landskap 2
19657 landskapen 1
19658 landskapet 1
19659 landsman 2
19660 landsmaninnor 2
19661 landsmän 6
19662 landsmäns 1
19663 landsspecifika 1
19664 landstiger 1
19665 landsväg 3
19666 landsändar 1
19667 landsätta 1
19668 landsättas 1
19669 landvinningar 4
19670 lansera 3
19671 lanserade 1
19672 lanserades 1
19673 lanserandet 1
19674 lanserar 1
19675 lanserat 1
19676 lansering 1
19677 lantbrukarna 1
19678 lantbruket 1
19679 lantbrukssamhälle 1
19680 lantdjur 1
19681 lantliga 1
19682 lappa 1
19683 lapptäcke 1
19684 lappverk 2
19685 larm 3
19686 larmrapporter 2
19687 larmsignal 2
19688 larver 1
19689 last 6
19690 lasta 2
19691 lastas 1
19692 lastat 1
19693 lastbil 5
19694 lastbilar 6
19695 lastbilarna 2
19696 lastbilsförare 1
19697 lastbilskontroll 1
19698 lastbilsparken 1
19699 lastbilsstänkskärmar 1
19700 lastbilsägare 1
19701 lastbilsägarna 1
19702 lasten 5
19703 lastens 2
19704 lasternas 1
19705 lastning 1
19706 lastområde 1
19707 lastrester 4
19708 lastrum 1
19709 lastångare 1
19710 latent 1
19711 latinamerikanska 1
19712 latituder 2
19713 latmansgöra 1
19714 lava 1
19715 law 2
19716 lax 7
19717 laxanemi 5
19718 laxanläggningar 1
19719 laxar 1
19720 laxen 2
19721 laxens 1
19722 laxindustrin 1
19723 laxodlare 1
19724 laxodlingar 1
19725 laxodlingsindustrin 1
19726 laxodlingssektorn 2
19727 laxrosa 1
19728 laxsektorn 1
19729 layout 6
19730 layouten 4
19731 le 6
19732 leasa 1
19733 led 4
19734 leda 121
19735 ledamot 99
19736 ledamoten 59
19737 ledamotens 6
19738 ledamotsstadga 1
19739 ledamotsstadgan 1
19740 ledamöter 157
19741 ledamöterna 58
19742 ledamöternas 8
19743 ledamöters 2
19744 ledande 15
19745 ledardjuren 1
19746 ledare 23
19747 ledaren 3
19748 ledarens 1
19749 ledares 1
19750 ledarförmåga 1
19751 ledarna 10
19752 ledarposition 1
19753 ledarskap 4
19754 ledarskapet 1
19755 ledas 2
19756 ledd 1
19757 ledda 2
19758 ledde 22
19759 leder 87
19760 ledet 3
19761 lediga 1
19762 ledmotiv 1
19763 ledning 16
19764 ledningar 1
19765 ledningen 14
19766 ledningscentralen 1
19767 ledningsförmågan 1
19768 ledningsmässiga 1
19769 ledningsnivåer 1
19770 ledningssätt 2
19771 ledningssättet 1
19772 ledningsutövning 1
19773 leds 2
19774 ledsaga 2
19775 ledsen 8
19776 ledstjärna 2
19777 ledstjärnan 1
19778 ledtrådar 1
19779 leende 17
19780 leendet 2
19781 legal 7
19782 legala 7
19783 legale 2
19784 legalisera 1
19785 legaliserade 1
19786 legalitet 4
19787 legaliteten 2
19788 legalitetsprincip 2
19789 legalt 9
19790 legat 5
19791 lege 1
19792 legionärerna 1
19793 legitim 3
19794 legitima 12
19795 legitimera 2
19796 legitimerar 2
19797 legitimeras 2
19798 legitimering 3
19799 legitimitet 10
19800 legitimiteten 3
19801 legitimt 1
19802 lejda 1
19803 lejer 1
19804 leka 1
19805 lekarna 1
19806 lekbeståndens 1
19807 lekboll 1
19808 leker 3
19809 lekfullt 1
19810 lekområde 1
19811 lekplats 1
19812 leksaker 2
19813 lekt 1
19814 lekte 4
19815 lektion 1
19816 lektioner 3
19817 lem 1
19818 lemlästande 1
19819 lemlästar 1
19820 lenande 1
19821 leninism 1
19822 ler 1
19823 lera 1
19824 leran 1
19825 lerhydda 1
19826 lerkärlen 1
19827 lerväggarna 1
19828 les 1
19829 leta 6
19830 letade 3
19831 letar 2
19832 lett 35
19833 leva 49
19834 levande 19
19835 levantinskt 1
19836 levat 1
19837 levde 6
19838 levebröd 5
19839 level 1
19840 lever 58
19841 leverans 1
19842 leverantör 1
19843 leverantörer 3
19844 leverantörskedjor 1
19845 leverar 1
19846 leverera 8
19847 levererar 2
19848 levereras 2
19849 levererat 3
19850 levnads- 1
19851 levnadsbetingelser 1
19852 levnadsglada 1
19853 levnadsnivå 1
19854 levnadsnivåer 1
19855 levnadsstandard 4
19856 levnadsstandarden 2
19857 levnadssätt 3
19858 levnadssättet 1
19859 levnadsvillkor 3
19860 levnadsvillkoren 1
19861 levt 3
19862 liaison 1
19863 libanesiska 1
19864 liberal 6
19865 liberala 56
19866 liberaldemokrater 1
19867 liberalen 1
19868 liberaler 3
19869 liberalerna 3
19870 liberalernas 1
19871 liberalisera 3
19872 liberalisering 4
19873 liberaliseringen 4
19874 liberalism 2
19875 liberalismen 2
19876 licens 1
19877 licenser 4
19878 licensfil 1
19879 licensiera 1
19880 licensinnehavarna 1
19881 licenspaketfil 1
19882 lida 6
19883 lidande 9
19884 lidanden 2
19885 lidandes 1
19886 lidandet 2
19887 lidelsefull 2
19888 lidelsefulla 4
19889 lider 21
19890 lidit 11
19891 lift 1
19892 liftare 1
19893 lifting 2
19894 liga 1
19895 ligga 34
19896 liggande 2
19897 ligger 179
19898 liggtidskostnaden 1
19899 lik 7
19900 lika 183
19901 likabehandling 1
19902 likaberättigad 1
19903 likadan 3
19904 likadana 3
19905 likadant 4
19906 likaledes 3
19907 likalydande 1
19908 likar 2
19909 likartad 1
19910 likartade 2
19911 likartat 1
19912 likaså 13
19913 likaväl 4
19914 likbleka 1
19915 likgiltig 2
19916 likgiltiga 3
19917 likgiltighet 2
19918 likgiltigheten 2
19919 likgiltigt 1
19920 likhet 33
19921 likheter 1
19922 likna 5
19923 liknade 7
19924 liknande 45
19925 liknar 12
19926 liknas 1
19927 liknat 1
19928 likriktade 4
19929 likriktande 1
19930 likriktas 1
19931 likriktning 2
19932 likriktningen 1
19933 liksidig 1
19934 liksom 157
19935 likstank 1
19936 likställa 3
19937 likställas 2
19938 likställda 2
19939 likställdes 1
19940 likställdhet 1
19941 likt 11
19942 likvida 2
19943 likväl 10
19944 likvärdig 4
19945 likvärdiga 8
19946 likvärdighet 1
19947 likvärdigt 1
19948 lila 1
19949 lilla 22
19950 lille 6
19951 lillfinger 2
19952 linan 1
19953 linbana 1
19954 linda 2
19955 lindra 4
19956 lindrande 1
19957 lindras 1
19958 lingua 1
19959 lingula 1
19960 lingvistiska 1
19961 linjal 1
19962 linje 34
19963 linjen 29
19964 linjer 5
19965 linjerna 4
19966 linjära 1
19967 linne 1
19968 linorna 1
19969 linsen 1
19970 lire 4
19971 lisa 1
19972 lista 13
19973 listan 13
19974 listigt 3
19975 listor 4
19976 listorna 2
19977 lita 6
19978 litade 2
19979 litar 9
19980 lite 28
19981 liten 63
19982 liter 1
19983 litet 145
19984 litteratur 6
19985 litteraturen 3
19986 litteraturförteckning 1
19987 litteraturförteckningen 1
19988 litterära 2
19989 liv 74
19990 livboj 1
19991 liverpoolskt 1
19992 livet 42
19993 livets 3
19994 livgardistuniform 1
19995 livlig 2
19996 livliga 5
19997 livligt 1
19998 livlina 2
19999 livnära 2
20000 livs 2
20001 livsbehov 2
20002 livsbesparingar 1
20003 livsbetingelserna 1
20004 livscykel 3
20005 livsdugliga 2
20006 livsförutsättningarna 1
20007 livshållning 1
20008 livskraft 2
20009 livskraften 1
20010 livskraftig 1
20011 livskraftiga 1
20012 livskvalitet 14
20013 livskvaliteten 9
20014 livskvalitén 2
20015 livslängden 1
20016 livslånga 1
20017 livslångt 9
20018 livsmedel 28
20019 livsmedels- 1
20020 livsmedelsbrist 2
20021 livsmedelsexport 1
20022 livsmedelsfrågor 1
20023 livsmedelsfrågorna 1
20024 livsmedelsföreskrifter 1
20025 livsmedelsföretagen 1
20026 livsmedelsförsörjningen 1
20027 livsmedelshanterares 1
20028 livsmedelshjälp 2
20029 livsmedelsindustrier 1
20030 livsmedelsindustrin 1
20031 livsmedelskedja 1
20032 livsmedelskedjan 2
20033 livsmedelskonsumtion 1
20034 livsmedelskontroll 2
20035 livsmedelskris 2
20036 livsmedelskriserna 1
20037 livsmedelskvalitet 3
20038 livsmedelslagstiftning 7
20039 livsmedelsmyndighet 8
20040 livsmedelsmyndigheten 4
20041 livsmedelsmyndighetens 1
20042 livsmedelsnyheterna 1
20043 livsmedelsområdet 1
20044 livsmedelsprodukter 1
20045 livsmedelsproduktion 1
20046 livsmedelsproduktionen 2
20047 livsmedelsproduktionskedjan 1
20048 livsmedelsprogram 1
20049 livsmedelssektorn 3
20050 livsmedelsstandarder 1
20051 livsmedelsstöd 1
20052 livsmedelssäkerhet 38
20053 livsmedelssäkerheten 7
20054 livsmedelssäkerhetens 1
20055 livsmedelssäkerhetsenheter 3
20056 livsmedelssäkerhetslagstiftningen 1
20057 livsmedelssäkerhetsmyndigheten 6
20058 livsmedelssäkerhetsmyndigheter 1
20059 livsmedelssäkerhetsområdet 1
20060 livsmedelssäkerhetssystem 1
20061 livsmedelstillverkningen 1
20062 livsmiljö 2
20063 livsmiljöer 6
20064 livsmiljöerna 1
20065 livsmiljön 1
20066 livsnödvändigt 1
20067 livspartner 1
20068 livsstil 1
20069 livstid 2
20070 livsuppehållande 1
20071 livsviktig 2
20072 livsviktigt 1
20073 livsvillkor 4
20074 livsyta 1
20075 livvakt 1
20076 ljud 6
20077 ljuda 1
20078 ljuder 1
20079 ljudet 3
20080 ljudlig 1
20081 ljudligt 1
20082 ljudlöst 1
20083 ljudupptagningar 6
20084 ljudupptagningar(11221/1999 1
20085 ljuga 2
20086 ljuger 1
20087 ljungeld 1
20088 ljus 18
20089 ljusa 4
20090 ljusan 1
20091 ljusare 2
20092 ljusblå 1
20093 ljusen 2
20094 ljuset 34
20095 ljushårig 1
20096 ljuskretsen 1
20097 ljuslagd 1
20098 ljuspunkter 1
20099 ljusrött 1
20100 ljussken 1
20101 ljusstråle 1
20102 ljustrafik 1
20103 ljusår 2
20104 ljuv 1
20105 ljuva 2
20106 ljuvlig 1
20107 ljuvliga 1
20108 ljuvligt 1
20109 lo 1
20110 lobby 1
20111 lobbyarbete 1
20112 lobbyarbetet 1
20113 lobbyföretag 1
20114 lobbygrupper 1
20115 lobbygrupperna 1
20116 lobbyintressen 1
20117 lobbymaskin 1
20118 lobbyverksamhet 3
20119 loca 1
20120 locka 4
20121 lockande 1
20122 lockar 1
20123 lockas 1
20124 lockats 1
20125 lockelse 2
20126 lockiga 1
20127 lockigt 2
20128 lodrät 1
20129 log 4
20130 logik 9
20131 logiken 5
20132 logisk 1
20133 logiska 4
20134 logiskt 13
20135 logistik 2
20136 logistiken 1
20137 logistikorganisation 1
20138 logistikstöd 1
20139 loj 1
20140 loja 1
20141 lojal 2
20142 lojalisterna 4
20143 lojalitet 1
20144 lojaliteten 1
20145 lojalt 3
20146 lojt 2
20147 lokal 27
20148 lokala 143
20149 lokalbefolkningen 2
20150 lokalen 1
20151 lokaler 4
20152 lokalerna 1
20153 lokaliseras 1
20154 lokalisering 2
20155 lokaliseringen 1
20156 lokaliseringsproblem 1
20157 lokalpatriotiska 1
20158 lokalpolis 1
20159 lokalsamhället 1
20160 lokalsamhällets 1
20161 lokalskatt 1
20162 lokalt 12
20163 lokaltidningen 1
20164 lokaltåg 1
20165 londonområdet 1
20166 look 1
20167 loopar 1
20168 lopp 9
20169 loppet 2
20170 loss 6
20171 lossa 1
20172 lossna 1
20173 lossnat 1
20174 lossning 1
20175 lots 1
20176 lotsat 1
20177 lotsens 1
20178 lotsning 1
20179 lott 2
20180 lottade 4
20181 lotusblomma 1
20182 lov 12
20183 lova 6
20184 lovade 17
20185 lovande 5
20186 lovar 7
20187 lovat 14
20188 lovats 1
20189 lovord 2
20190 lovorda 4
20191 lovordar 2
20192 lovordats 1
20193 lovprisar 1
20194 lovvärd 2
20195 lovvärda 3
20196 lovvärt 1
20197 lovyttringar 1
20198 lucka 4
20199 luckor 6
20200 luckorna 1
20201 luckra 1
20202 luddiga 3
20203 luddighet 1
20204 luddigt 2
20205 luft 5
20206 luftbro 1
20207 luftburet 1
20208 luftburna 1
20209 luften 18
20210 luftfarkost 1
20211 luftfart 1
20212 luftföroreningar 1
20213 luftkvalitet 1
20214 luftområde 1
20215 lufträder 1
20216 luftslottsbetänkande 1
20217 luftströmmarna 1
20218 lufttransport- 1
20219 lufttransporter 1
20220 lufttransporterna 1
20221 lugg 1
20222 luggar 1
20223 luggslitna 1
20224 lugn 8
20225 lugna 11
20226 lugnade 3
20227 lugnande 2
20228 lugnar 3
20229 lugnare 1
20230 lugnas 1
20231 lugnt 4
20232 lukrativa 1
20233 lukt 1
20234 luktade 4
20235 luktar 1
20236 lukten 2
20237 lukter 1
20238 lumpsamlarverksamhet 1
20239 lunch 2
20240 lunchen 2
20241 luncher 1
20242 lunchtid 1
20243 lungor 1
20244 lur 1
20245 lura 1
20246 lurad 1
20247 lurande 1
20248 luras 3
20249 lurat 1
20250 luren 4
20251 lust 6
20252 lusten 1
20253 lustiga 3
20254 lustigare 1
20255 lustigt 1
20256 luta 2
20257 lutad 1
20258 lutade 9
20259 lutande 1
20260 lutar 1
20261 lutheranska 1
20262 lutning 1
20263 luxemburgare 1
20264 luxemburgska 1
20265 lycka 9
20266 lyckad 2
20267 lyckade 5
20268 lyckades 25
20269 lyckan 3
20270 lyckas 77
20271 lyckat 2
20272 lyckats 52
20273 lycklig 11
20274 lyckliga 4
20275 lyckligaste 1
20276 lyckligt 2
20277 lyckligtvis 6
20278 lyckojägare 1
20279 lyckosamt 2
20280 lyckönska 7
20281 lyckönskas 1
20282 lyckönskningar 5
20283 lyckönskningsmeddelande 1
20284 lyda 4
20285 lydelse 4
20286 lyder 15
20287 lydigt 1
20288 lydnad 1
20289 lyft 3
20290 lyfta 19
20291 lyftade 1
20292 lyftas 1
20293 lyfte 8
20294 lyfter 3
20295 lyftkraftsteori 1
20296 lyhörd 1
20297 lyhördhet 2
20298 lykta 1
20299 lyktornas 1
20300 lynchad 1
20301 lynchningsscener 1
20302 lyrisk 1
20303 lyriska 1
20304 lysa 4
20305 lysande 9
20306 lyser 3
20307 lyssna 32
20308 lyssnade 14
20309 lyssnande 1
20310 lyssnar 13
20311 lyssnat 20
20312 lyssningsläge 1
20313 lyst 1
20314 lyste 2
20315 lyxproblem 1
20316 läck 1
20317 läcka 2
20318 läckage 2
20319 läckan 1
20320 läckande 2
20321 läcker 4
20322 läckor 2
20323 läckt 4
20324 läckte 3
20325 läder 1
20326 läderpåse 1
20327 läge 28
20328 lägen 1
20329 lägena 1
20330 lägenhet 1
20331 lägenheten 7
20332 läger 2
20333 lägesbedömningar 1
20334 lägesrapport 2
20335 läget 24
20336 lägg 2
20337 lägga 204
20338 läggas 22
20339 lägger 76
20340 läggning 2
20341 läggs 45
20342 läglig 1
20343 lägliga 1
20344 lägligt 4
20345 lägre 26
20346 lägret 1
20347 lägst 2
20348 lägsta 7
20349 läkare 6
20350 läkarjobb 1
20351 läkarkontroller 2
20352 läkartjänst 1
20353 läkemedel 4
20354 läkemedelsindustrin 1
20355 läktarna 1
20356 lämna 68
20357 lämnad 2
20358 lämnade 14
20359 lämnades 3
20360 lämnar 30
20361 lämnas 17
20362 lämnat 25
20363 lämnats 9
20364 lämningarna 1
20365 lämpa 1
20366 lämpade 3
20367 lämpar 2
20368 lämplig 27
20369 lämpliga 38
20370 lämpligare 4
20371 lämpligast 1
20372 lämpligaste 3
20373 lämpligen 1
20374 lämplighet 2
20375 lämpligheten 1
20376 lämplighetsprov 1
20377 lämpligt 66
20378 län 2
20379 länder 361
20380 länderna 135
20381 ländernas 18
20382 länders 14
20383 ländskynken 1
20384 längd 3
20385 längden 3
20386 länge 124
20387 längesedan 2
20388 längre 204
20389 längs 26
20390 längst 5
20391 längsta 1
20392 längtan 2
20393 längtar 2
20394 länk 10
20395 länka 3
20396 länkad 2
20397 länkade 1
20398 länken 1
20399 läppar 4
20400 läpparna 1
20401 läpparnas 1
20402 läppstift 1
20403 lär 7
20404 lära 34
20405 lärande 11
20406 lärandet 2
20407 lärare 4
20408 läraren 1
20409 lärarna 3
20410 läras 1
20411 lärd 1
20412 lärda 1
20413 lärde 4
20414 lärdom 13
20415 lärdomar 4
20416 läroanstalter 1
20417 läroplanen 1
20418 lärorikt 1
20419 lärosatser 1
20420 lärs 1
20421 lärt 12
20422 lärts 1
20423 läs 3
20424 läsa 11
20425 läsas 1
20426 läsbar 1
20427 läsbara 1
20428 läsbarare 1
20429 läser 23
20430 läsfrämjande 1
20431 läskunniga 1
20432 läskunnigheten 1
20433 läsningen 1
20434 läst 11
20435 läste 13
20436 lät 14
20437 lätt 52
20438 lätta 7
20439 lättad 1
20440 lättade 1
20441 lättar 2
20442 lättare 38
20443 lättast 2
20444 lättaste 1
20445 lättflytande 1
20446 lättförståelig 1
20447 lättförståeligt 1
20448 lätthet 1
20449 lättillgänglig 1
20450 lättillgängliga 1
20451 lättläst 1
20452 lättnad 3
20453 lättnader 3
20454 lättrogenhet 1
20455 lättsinnig 1
20456 lättsinnigt 1
20457 lättviktsfordon 1
20458 lättviktsmetoder 1
20459 lättvättat 1
20460 läxa 4
20461 läxan 3
20462 läxat 1
20463 läxor 4
20464 lådfacks 1
20465 lådor 1
20466 lådorna 1
20467 låg 60
20468 låga 24
20469 låginkomsttagare 2
20470 låglönestrategierna 1
20471 lågorna 1
20472 lågt 9
20473 lån 3
20474 låna 1
20475 lånade 1
20476 lånat 1
20477 lånats 1
20478 lång 109
20479 lång- 1
20480 långa 52
20481 långdragen 2
20482 långdragna 1
20483 långfenad 1
20484 långfingret 1
20485 långfristig 1
20486 långfärdsbussar 1
20487 långrandig 2
20488 långrandigt 1
20489 långsam 1
20490 långsamhet 1
20491 långsamheten 1
20492 långsamma 6
20493 långsammare 3
20494 långsamt 20
20495 långsiktig 5
20496 långsiktiga 18
20497 långsiktighet 1
20498 långsiktigt 9
20499 långt 113
20500 långtgående 14
20501 långtids- 1
20502 långtidsarbetslösa 4
20503 långtidsarbetslöshet 5
20504 långtidsarbetslösheten 1
20505 långtifrån 3
20506 långtradare 2
20507 långvariga 8
20508 långvarigt 4
20509 låsa 4
20510 låser 1
20511 låset 1
20512 låsningarna 1
20513 låsningen 1
20514 låst 2
20515 låsta 1
20516 låsts 1
20517 låt 47
20518 låta 102
20519 låter 32
20520 låtit 6
20521 låtsad 1
20522 låtsades 1
20523 låtsas 9
20524 löddrade 1
20525 löfte 14
20526 löften 21
20527 löftena 1
20528 löftesrika 1
20529 löftesrikt 1
20530 löftet 4
20531 lögn 1
20532 lögnen 1
20533 lögner 2
20534 löjeväckande 4
20535 löjliga 1
20536 lökar 1
20537 lökformade 2
20538 lökmodell 1
20539 lömsk 1
20540 lömskt 1
20541 lön 8
20542 löna 2
20543 lönar 1
20544 löne- 3
20545 lönearbetsrättigheter 1
20546 lönebesked 2
20547 löneeffektivitet 1
20548 löneförhållandena 1
20549 lönehöjningarna 1
20550 lönemässigt 1
20551 lönen 2
20552 lönepaketet 1
20553 lönepolitik 3
20554 löner 8
20555 lönerna 2
20556 lönetak 1
20557 löneökningar 1
20558 löneökningspolitik 1
20559 lönsam 3
20560 lönsamhet 2
20561 lönsamhets- 1
20562 lönsamhetstänkande 1
20563 lönsamma 6
20564 lönsamt 2
20565 lönt 2
20566 löntagare 2
20567 löntagarna 6
20568 löpa 4
20569 löpande 11
20570 löpeld 1
20571 löper 12
20572 löpt 6
20573 löpte 5
20574 lördag 1
20575 lördagskvällar 1
20576 lös 5
20577 lösa 103
20578 lösare 1
20579 lösas 16
20580 löser 9
20581 löses 2
20582 lösesumma 1
20583 lösgör 1
20584 lösning 109
20585 lösningar 51
20586 lösningarna 1
20587 lösningen 23
20588 lösningsförslag 1
20589 lösnäsa 1
20590 lösryckt 1
20591 löst 10
20592 lösta 5
20593 löste 2
20594 löstes 3
20595 lösts 8
20596 löv 1
20597 lövskogarna 1
20598 m 1
20599 m.fl. 3
20600 m.m. 5
20601 m3 2
20602 mader 1
20603 maffia 1
20604 maffian 1
20605 maffians 1
20606 maffior 1
20607 magasin 3
20608 magasinerade 2
20609 mage 1
20610 magen 4
20611 mager 5
20612 magi 3
20613 magisk 1
20614 magiska 1
20615 magiskt 1
20616 magnet 1
20617 magnifik 1
20618 magnifika 1
20619 magnitud 1
20620 magra 1
20621 magrare 1
20622 magstarkt 1
20623 mainstraming 1
20624 mainstreaming 18
20625 mainstreaming-program 1
20626 maj 23
20627 majestätiskt 1
20628 majoritet 54
20629 majoriteten 19
20630 majoriteter 1
20631 majoritetsbeslut 4
20632 majoritetsbeslutet 1
20633 majoritetsgrupp 1
20634 majoritetsomröstningar 1
20635 majoritetsröstning 1
20636 majoritetsuppfattning 1
20637 majoritetsuppfattningen 1
20638 makabert 1
20639 makade 1
20640 makarna 2
20641 make 2
20642 makedonierna 3
20643 makedonisk 1
20644 makedoniska 7
20645 makedoniskt 1
20646 maken 1
20647 makroekonomin 1
20648 makroekonomisk 5
20649 makroekonomiska 17
20650 makroekonomiskt 3
20651 makrofinansiellt 1
20652 makropolitik 1
20653 makt 40
20654 maktambitioner 1
20655 maktbalans 1
20656 maktbalansen 1
20657 maktbefogenhet 3
20658 maktbefogenheter 2
20659 maktberusning 1
20660 maktcentrumen 1
20661 maktdelningen 1
20662 maktdikterade 1
20663 makten 23
20664 maktens 2
20665 makter 2
20666 makterna 1
20667 maktfaktor 2
20668 maktförlusten 1
20669 makthavare 2
20670 makthavarna 2
20671 maktkoncentration 2
20672 maktkoncentrationen 1
20673 maktkoncentrationer 1
20674 maktlös 4
20675 maktlösa 1
20676 maktlöshet 3
20677 maktlöst 1
20678 maktmedel 3
20679 maktmedlen 1
20680 maktmissbruk 3
20681 maktpolitiska 1
20682 maktpositionen 1
20683 maktpositioner 2
20684 maktstrukturer 1
20685 maktövertagande 1
20686 mal 1
20687 malaria 1
20688 malariamyggan 1
20689 maldes 1
20690 mall 3
20691 malplacerade 1
20692 malt 1
20693 maltesarna 1
20694 malteserna 1
20695 maltesisk 3
20696 maltesiska 2
20697 maltwhisky 1
20698 maltwhiskyproducerande 1
20699 mamma 6
20700 man 1871
20701 mana 2
20702 manad 1
20703 manade 1
20704 management 1
20705 managementnivå 1
20706 manar 4
20707 manas 1
20708 manat 1
20709 mandat 18
20710 mandaten 1
20711 mandatet 4
20712 mandatperiod 15
20713 mandatperioden 10
20714 mandatperiodens 2
20715 maner 1
20716 mangoträden 1
20717 mangoträdens 1
20718 mangroveträden 1
20719 manifestationen 1
20720 manifestationer 1
20721 manifestationerna 1
20722 manifesterar 1
20723 maning 2
20724 manipulation 2
20725 manipulerad 1
20726 manlig 2
20727 manliga 10
20728 manligt 1
20729 manna 1
20730 mannen 18
20731 mannens 2
20732 mans 1
20733 manschettknappar 1
20734 mantra 1
20735 mantran 1
20736 mantrat 1
20737 manuellt 1
20738 manuskriptet 1
20739 manér 1
20740 manöver 2
20741 manövern 1
20742 manövrer 1
20743 manövrerade 1
20744 mapp 1
20745 mapparna 2
20746 mappen 2
20747 maratonlångt 1
20748 mardrömmar 3
20749 mardrömslik 1
20750 marginal 3
20751 marginalen 3
20752 marginaler 3
20753 marginalerna 1
20754 marginalisera 3
20755 marginaliserade 5
20756 marginaliserats 1
20757 marginalisering 2
20758 marginellt 2
20759 marin 2
20760 marina 18
20761 marionett 1
20762 maritima 2
20763 maritimt 2
20764 mark 13
20765 markant 4
20766 markanta 1
20767 markanvändning 1
20768 marken 12
20769 markens 1
20770 markera 2
20771 markerad 1
20772 markerade 1
20773 markerades 1
20774 markerar 9
20775 markeras 2
20776 markerat 2
20777 markering 2
20778 market 1
20779 marknad 50
20780 marknaden 190
20781 marknadens 26
20782 marknader 21
20783 marknaderna 18
20784 marknadernas 7
20785 marknadsaktören 1
20786 marknadsaktörerna 1
20787 marknadsaktörernas 1
20788 marknadsandel 2
20789 marknadsandelar 8
20790 marknadsdominans 1
20791 marknadsekonomi 13
20792 marknadsekonomin 8
20793 marknadsekonomins 2
20794 marknadsekonomiska 3
20795 marknadsföring 2
20796 marknadsföringskoncept 1
20797 marknadsinstrumentet 1
20798 marknadskrafter 1
20799 marknadskrafterna 1
20800 marknadslagarna 1
20801 marknadsliberalism 1
20802 marknadsmöjlighet 1
20803 marknadsorganisation 1
20804 marknadsorganisationen 1
20805 marknadspriser 2
20806 marknadsproblem 2
20807 marknadsprodukt 1
20808 marknadssituation 1
20809 marknadstillträde 4
20810 marktrupper 1
20811 marmorbyggnad 1
20812 marmortrappan 1
20813 marockanska 4
20814 marokäng 1
20815 mars 55
20816 marschera 1
20817 marscherande 1
20818 marscherar 1
20819 marshmallow 1
20820 marshmallow-klunsar 1
20821 marshmallowen 1
20822 marshmallows 1
20823 marskgräs 1
20824 marskgräset 2
20825 martinis 1
20826 mask 1
20827 masker 1
20828 maskerad 1
20829 maskin 3
20830 maskinellt 1
20831 maskinen 1
20832 maskiner 1
20833 maskineri 2
20834 maskineriet 2
20835 maskinist 1
20836 maskinistexamen 1
20837 maskinrummen 1
20838 maskinrummet 1
20839 maskinskada 1
20840 maskopi 1
20841 maskstungna 1
20842 masochister 1
20843 masochistisk 1
20844 masochistiska 1
20845 massa 11
20846 massakerplatserna 1
20847 massakrera 1
20848 massakrerade 1
20849 massakrerna 1
20850 massan 1
20851 massans 1
20852 massarbetslöshet 1
20853 massarbetslösheten 2
20854 massavgång 1
20855 massiv 3
20856 massiva 7
20857 massivt 2
20858 massmedia 4
20859 massmedias 2
20860 massrörelse 1
20861 masten 1
20862 masterna 1
20863 mastodont 1
20864 mat 11
20865 mata 1
20866 match 1
20867 matcha 2
20868 matchande 1
20869 matchar 2
20870 matdags 1
20871 matematiker 1
20872 matematisk 1
20873 matematiska 1
20874 maten 3
20875 material 28
20876 materialanskaffning 1
20877 materialen 1
20878 materialet 3
20879 materiell 1
20880 materiella 2
20881 materiellt 2
20882 matlagning 1
20883 matnyttiga 1
20884 matpaket 2
20885 matpensioner 1
20886 matrester 1
20887 matroserna 1
20888 matsal 1
20889 matsalen 1
20890 matsedeln 1
20891 matsedlarna 1
20892 matt 1
20893 matta 1
20894 mattan 2
20895 mattorna 1
20896 maxbeloppen 1
20897 maximal 7
20898 maximala 3
20899 maximalt 7
20900 maximera 4
20901 maximerar 1
20902 maximistraffet 1
20903 maxstraffet 1
20904 maxvikter 1
20905 med 5080
20906 medaljbehängda 1
20907 medan 107
20908 medansvar 3
20909 medarbetare 7
20910 medbeslutande 14
20911 medbeslutandeförfarande 3
20912 medbeslutandeförfarandet 11
20913 medbeslutanderätt 3
20914 medbeslutandet 3
20915 medborgardebatt 1
20916 medborgardebatter 1
20917 medborgardemonstration 1
20918 medborgare 142
20919 medborgaren 21
20920 medborgaren-konsumenten 1
20921 medborgarens 1
20922 medborgares 18
20923 medborgarna 170
20924 medborgarnas 59
20925 medborgarrätt 1
20926 medborgarrörelser 1
20927 medborgarsamhället 2
20928 medborgarskap 6
20929 medborgarskapet 4
20930 medborgarskapsbegrepp 1
20931 medborgarskapsregleringen 1
20932 medborgarstadga 1
20933 medborgartanken 1
20934 medborgarvärde 1
20935 medborgerlig 1
20936 medborgerliga 21
20937 medborgerligt 2
20938 medbroders 1
20939 medbrottslighet 1
20940 medbrottslingar 1
20941 meddela 25
20942 meddelade 7
20943 meddelades 1
20944 meddelande 89
20945 meddelanden 12
20946 meddelandeskyldigheten 1
20947 meddelandet 34
20948 meddelandetexten 1
20949 meddelar 7
20950 meddelat 5
20951 medel 165
20952 medel- 1
20953 medelklass 3
20954 medellängd 1
20955 medellång 13
20956 medelmåttan 1
20957 medelmåttiga 1
20958 medelpunkt 2
20959 medelst 1
20960 medelstor 3
20961 medelstora 72
20962 medelstort 1
20963 medeltida 3
20964 medeltiden 1
20965 medelvärden 1
20966 medelålder 1
20967 medelåldern 1
20968 medelålders 1
20969 medfarna 1
20970 medfinansierade 1
20971 medfinansieras 1
20972 medfinansiering 1
20973 medfinansieringen 1
20974 medföljde 1
20975 medför 43
20976 medföra 17
20977 medförde 3
20978 medföredragande 2
20979 medfört 5
20980 medgav 2
20981 medge 7
20982 medger 24
20983 medges 9
20984 medgett 1
20985 medgivande 2
20986 medgivits 2
20987 medgörliga 1
20988 medgörlighet 1
20989 medhjälpare 1
20990 media 11
20991 mediaföretagen 1
20992 medial 1
20993 mediatäckningen 1
20994 medicin 2
20995 mediciner 1
20996 medicinsk 3
20997 medicinska 1
20998 medie- 1
20999 medier 7
21000 medierna 4
21001 mediernas 3
21002 medinflytande 2
21003 meditera 1
21004 medkänsla 9
21005 medla 2
21006 medlare 1
21007 medlaren 1
21008 medlem 23
21009 medlemmar 41
21010 medlemmarna 2
21011 medlemmars 1
21012 medlemsavgifter 1
21013 medlemskandidaterna 1
21014 medlemskap 23
21015 medlemskapet 1
21016 medlemskapsförhandlingarna 4
21017 medlemskapsprocessen 2
21018 medlemskapsrättigheter 1
21019 medlemskapsstöden 1
21020 medlemskapsåtgärder 1
21021 medlemsland 12
21022 medlemslandet 3
21023 medlemslands 1
21024 medlemsländer 21
21025 medlemsländerna 38
21026 medlemsländernas 12
21027 medlemsländers 2
21028 medlemsregeringarnas 1
21029 medlemsstarter 1
21030 medlemsstat 88
21031 medlemsstaten 15
21032 medlemsstatens 3
21033 medlemsstater 196
21034 medlemsstaterna 329
21035 medlemsstaterna- 1
21036 medlemsstaternas 90
21037 medlemsstaters 9
21038 medlemsstats 13
21039 medlemsstatsnivå 7
21040 medlemsstatsrapport 1
21041 medlen 20
21042 medlet 2
21043 medlidande 2
21044 medling 1
21045 medlingsförfarande 3
21046 medlingsförsök 1
21047 medlingsförsöken 1
21048 medlingsprocess 1
21049 medmänniskors 1
21050 medmänskliga 1
21051 medmänsklighet 2
21052 medskyldiga 2
21053 medspelarna 1
21054 medsvuren 1
21055 medverka 17
21056 medverkade 1
21057 medverkan 12
21058 medverkar 9
21059 medverkat 4
21060 medvetande 8
21061 medvetandehöjande 1
21062 medvetandenivå 1
21063 medvetandet 1
21064 medveten 46
21065 medvetenhet 7
21066 medvetenheten 1
21067 medvetet 12
21068 medvetna 59
21069 megaprojekt 1
21070 mej 1
21071 mejeriindustrin 1
21072 meka 1
21073 mekanik 1
21074 mekanisk 2
21075 mekaniska 3
21076 mekaniskt 3
21077 mekanism 5
21078 mekanismen 1
21079 mekanismer 18
21080 mekanismerna 7
21081 mekanistiska 1
21082 mellan 721
21083 mellanfolklig 1
21084 mellanlagras 1
21085 mellanlagringar 1
21086 mellanled 2
21087 mellanliggande 5
21088 mellannivå 1
21089 mellanrum 1
21090 mellanskillnaden 1
21091 mellanstadiet 1
21092 mellanstatlig 5
21093 mellanstatliga 2
21094 mellanstatligt 6
21095 mellanstora 2
21096 mellanting 1
21097 mellanvägg 1
21098 mellanöstern 1
21099 membre 2
21100 memoarer 1
21101 men 1306
21102 mena 1
21103 menade 12
21104 menar 69
21105 menas 3
21106 mening 91
21107 meningar 3
21108 meningarna 1
21109 meningen 16
21110 meningsfull 4
21111 meningsfulla 3
21112 meningsfullt 14
21113 meningslös 4
21114 meningslösa 2
21115 meningslöst 7
21116 meningsskiljaktigheter 8
21117 meningsskiljaktigheterna 1
21118 menligt 1
21119 mentalitet 1
21120 mentaliteten 5
21121 mentalsjuk 1
21122 meny 1
21123 mer 602
21124 mera 60
21125 merger 1
21126 meriter 4
21127 meritokrati 1
21128 merkostnaden 1
21129 merparten 1
21130 mervärde 10
21131 mervärdesskattesats 1
21132 mervärdesstruktur 1
21133 mervärdet 1
21134 mesanmasten 1
21135 mest 146
21136 mesta 11
21137 mestadels 2
21138 metaforen 1
21139 metafysiskt 1
21140 metall 1
21141 metaller 3
21142 metallindustrin 1
21143 metalliska 1
21144 meter 2
21145 metersystemet 1
21146 metervis 1
21147 metod 29
21148 metoden 8
21149 metoder 36
21150 metoderna 5
21151 metodik 1
21152 metodiken 3
21153 metodikens 1
21154 metodikändringar 1
21155 metodiskt 4
21156 metodutveckling 1
21157 middag 4
21158 middagen 6
21159 middagsbjudningen 1
21160 middagsbord 1
21161 middagshetta 1
21162 midja 1
21163 midjan 2
21164 midnatt 2
21165 mig 752
21166 migration 2
21167 migrationen 2
21168 migrationsrörelser 1
21169 migrationsströmmar 2
21170 migrationsströmmen 1
21171 mikrober 1
21172 mikroföretag 2
21173 mikrokrediter 2
21174 mikroprojekt 1
21175 mikrostater 1
21176 mikrostaterna 1
21177 mild 1
21178 mildare 1
21179 mildaste 1
21180 mildra 8
21181 mildrande 1
21182 mildras 1
21183 milen 1
21184 milis 2
21185 militariserade 1
21186 militarisering 2
21187 militarismen 1
21188 militär 19
21189 militära 52
21190 militäraktion 1
21191 militäraktioner 1
21192 militärer 2
21193 militärerna 1
21194 militärindustri 1
21195 militärinsats 1
21196 militärinsatserna 1
21197 militärkupp 1
21198 militärläger 1
21199 militärpolitiken 1
21200 militärsamarbete 1
21201 militärstyrkorna 1
21202 militärstyrkornas 1
21203 militärt 4
21204 militäruniformer 1
21205 miljard 1
21206 miljarder 40
21207 miljon 10
21208 miljoner 176
21209 miljonerna 2
21210 miljontals 3
21211 miljö 98
21212 miljö- 7
21213 miljöanpassad 2
21214 miljöansvar 3
21215 miljöansvaret 2
21216 miljöansvariga 1
21217 miljöarbete 1
21218 miljöarbetet 3
21219 miljöaspekten 4
21220 miljöaspekter 1
21221 miljöaspekterna 5
21222 miljöavtal 1
21223 miljöbelastningen 1
21224 miljöberoendet 1
21225 miljöbeskattning 1
21226 miljöbeskattningen 1
21227 miljöbestämmelser 1
21228 miljöbestämmelserna 1
21229 miljöbovar 1
21230 miljöbovarna 1
21231 miljöbrott 1
21232 miljöbrottsmyndighet 1
21233 miljöcowboys 1
21234 miljödepartementet 1
21235 miljödimensionen 2
21236 miljödirektiv 3
21237 miljödirektiven 1
21238 miljödirektivet 1
21239 miljödirektoratet 1
21240 miljödogmatism 1
21241 miljöeffekter 1
21242 miljöer 5
21243 miljöexperter 1
21244 miljöfaktor 1
21245 miljöfarliga 1
21246 miljöfråga 1
21247 miljöfrågan 1
21248 miljöfrågor 11
21249 miljöfrågorna 3
21250 miljöförbättrande 1
21251 miljöförbättring 1
21252 miljöfördelar 1
21253 miljöförhållandena 1
21254 miljöförordningen 1
21255 miljöförstörande 1
21256 miljöförstörelse 2
21257 miljöförstöring 5
21258 miljöförstöringen 1
21259 miljöförsämring 1
21260 miljögrupper 1
21261 miljöhänsyn 10
21262 miljöhänsynen 1
21263 miljöinformation 1
21264 miljöinsatserna 1
21265 miljökastastrofen 1
21266 miljökatastrof 12
21267 miljökatastrofala 1
21268 miljökatastrofen 3
21269 miljökatastrofens 1
21270 miljökatastroferna 1
21271 miljökommissionär 1
21272 miljökommissionären 1
21273 miljökonferensen 1
21274 miljökonsekvensbedömning 2
21275 miljökonsekvensbeskrivning 1
21276 miljökonsekvenser 5
21277 miljökonsekvenserna 3
21278 miljökostnaderna 2
21279 miljökrav 6
21280 miljökraven 4
21281 miljökunskap 1
21282 miljökvaliteten 1
21283 miljölagstiftning 3
21284 miljölagstiftningen 2
21285 miljölagstiftningens 1
21286 miljömedvetandet 2
21287 miljömetoder 1
21288 miljöminister 3
21289 miljöministern 1
21290 miljöministrarna 1
21291 miljömyndigheterna 1
21292 miljömässig 2
21293 miljömässiga 18
21294 miljömässigt 5
21295 miljömål 5
21296 miljömålen 1
21297 miljömålsättningarna 1
21298 miljön 122
21299 miljönormer 2
21300 miljönormerna 2
21301 miljöns 3
21302 miljönätverk 1
21303 miljöområde 1
21304 miljöområden 2
21305 miljöområdet 13
21306 miljöorgan 1
21307 miljöorganisation 1
21308 miljöovänligt 1
21309 miljöpartist 1
21310 miljöpelaren 1
21311 miljöperspektiv 1
21312 miljöpolicyavtal 1
21313 miljöpolitik 7
21314 miljöpolitiken 7
21315 miljöpolitikens 1
21316 miljöpolitisk 1
21317 miljöpolitiska 2
21318 miljöpolitiskt 3
21319 miljöproblem 5
21320 miljöproblemen 3
21321 miljöprogram 1
21322 miljöprogrammen 1
21323 miljöprogrammering 1
21324 miljöprojekt 1
21325 miljöpåverkan 4
21326 miljöregelverket 1
21327 miljörelaterade 1
21328 miljöresultat 1
21329 miljörisker 1
21330 miljörådet 1
21331 miljörörelsen 3
21332 miljörörelsens 1
21333 miljörörelserna 1
21334 miljösektorerna 1
21335 miljösidan 1
21336 miljösituationen 1
21337 miljöskadliga 2
21338 miljöskador 2
21339 miljöskydd 16
21340 miljöskyddet 5
21341 miljöskyddets 1
21342 miljöskyddsbehoven 1
21343 miljöskyddsnivå 2
21344 miljöskyddsområdet 1
21345 miljöskyddspolitik 1
21346 miljöskyddsstöd 1
21347 miljöskäl 3
21348 miljöstudier 1
21349 miljöstöd 1
21350 miljösyften 1
21351 miljösynpunkt 8
21352 miljötragedi 1
21353 miljötvånget 1
21354 miljöuppgifter 2
21355 miljöutskottet 7
21356 miljövariabler 1
21357 miljövänlig 2
21358 miljövänliga 7
21359 miljövänligaste 1
21360 miljövänligt 4
21361 miljövärdena 2
21362 miljöövervakningsenhet 1
21363 milkshakes 1
21364 millenniefebern 1
21365 millenniefusioner 1
21366 millennieskifte 1
21367 millennieskiftet 2
21368 millenniet 4
21369 millennietal 1
21370 millenniets 1
21371 millennium 2
21372 millimeteranpassade 1
21373 milstolpar 1
21374 milstolpe 3
21375 min 479
21376 min. 1
21377 mina 207
21378 minamatasjukdomen 1
21379 mindervärdiga 1
21380 minderårig 1
21381 minderåriga 1
21382 mindes 3
21383 mindre 181
21384 mineraler 1
21385 miniatyr 2
21386 minimal 1
21387 minimala 1
21388 minimalistiska 1
21389 minimalistiskt 1
21390 minimera 6
21391 minimeras 1
21392 minimibelopp 1
21393 minimibestämmelser 2
21394 minimifinansiering 1
21395 minimigemenskapsprogram 1
21396 minimiinkomst 1
21397 minimiinnehållet 1
21398 minimiinsatser 1
21399 minimikalender 1
21400 minimikapital 1
21401 minimikontroll 1
21402 minimikrav 4
21403 minimikraven 1
21404 minimikvoter 1
21405 minimilängden 1
21406 minimilön 1
21407 minimilönen 1
21408 minimilöner 2
21409 miniminivå 2
21410 miniminivån 1
21411 miniminormer 5
21412 minimipensionerna 1
21413 minimiprogram 1
21414 minimiprogrammet 2
21415 minimireform 2
21416 minimireformer 1
21417 minimiregler 5
21418 minimireglerna 2
21419 minimirättigheterna 1
21420 minimis-notis 1
21421 minimiskatter 1
21422 minimistandarden 1
21423 minimistandarder 2
21424 minimitaket 1
21425 minimitarifferna 1
21426 minimiuppehälle 1
21427 minimivikt 1
21428 minimiåtgärder 1
21429 minimorum 1
21430 minimum 12
21431 minireform 1
21432 minister 17
21433 ministerier 1
21434 ministermöte 1
21435 ministermötet 3
21436 ministern 16
21437 ministernivå 1
21438 ministerns 1
21439 ministerpost 1
21440 ministerposter 2
21441 ministerpresidenten 3
21442 ministerråd 5
21443 ministerrådet 22
21444 ministerrådets 1
21445 ministerrådsmöte 1
21446 ministrar 16
21447 ministrarna 8
21448 ministrars 1
21449 mink 1
21450 minkpäls 1
21451 minnas 6
21452 minne 11
21453 minnen 2
21454 minnena 1
21455 minnens 1
21456 minnesbild 1
21457 minnesmärke 1
21458 minnesvärda 1
21459 minnet 9
21460 minns 20
21461 minore 1
21462 minoritet 16
21463 minoriteten 7
21464 minoritetens 1
21465 minoriteter 25
21466 minoriteterna 6
21467 minoriteternas 2
21468 minoriteters 2
21469 minoritetsbefolkningar 1
21470 minoritetsfientliga 1
21471 minoritetsgrupper 5
21472 minoritetspolitik 1
21473 minoritetspolitiken 1
21474 minoritetsregering 3
21475 minorna 1
21476 minpolitiken 1
21477 minröjning 1
21478 minsann 2
21479 minska 86
21480 minskad 13
21481 minskade 11
21482 minskades 2
21483 minskande 4
21484 minskar 26
21485 minskas 9
21486 minskat 17
21487 minskats 2
21488 minskning 37
21489 minskningar 3
21490 minskningen 8
21491 minst 97
21492 minsta 29
21493 minste 1
21494 minttabletter 1
21495 minus 3
21496 minusgrader 2
21497 minut 13
21498 minuten 2
21499 minuter 21
21500 minåtgärdsprogrammens 1
21501 mirakel 1
21502 mirakellösning 1
21503 mirakelmedel 1
21504 mirakulöst 1
21505 missa 2
21506 missade 2
21507 missat 4
21508 missbelåtenhet 1
21509 missbruk 14
21510 missbruka 1
21511 missbrukade 1
21512 missbrukades 1
21513 missbrukar 1
21514 missbrukas 1
21515 missbrukat 1
21516 missbruket 2
21517 missbruksprincipen 1
21518 missfall 1
21519 missfallen 2
21520 missfoster 1
21521 missförhållande 2
21522 missförhållandena 1
21523 missförhållandet 1
21524 missförstod 2
21525 missförstå 1
21526 missförstånd 7
21527 missförstår 1
21528 missförstås 1
21529 missgynna 2
21530 missgynnade 14
21531 missgynnas 1
21532 misshandel 3
21533 misshandlade 1
21534 misshandlar 1
21535 misshushållning 2
21536 mission 2
21537 missions 1
21538 missionären 1
21539 misskreditera 1
21540 misskrediterar 1
21541 misskötsel 7
21542 misskött 1
21543 misslyckad 1
21544 misslyckade 5
21545 misslyckades 5
21546 misslyckande 13
21547 misslyckanden 5
21548 misslyckandet 2
21549 misslyckas 14
21550 misslyckat 1
21551 misslyckats 9
21552 missnöjd 2
21553 missnöjda 1
21554 missnöje 4
21555 missta 1
21556 misstag 17
21557 misstagen 3
21558 misstaget 2
21559 misstankar 6
21560 misstanke 2
21561 misstar 3
21562 misstolkas 2
21563 misstro 5
21564 misstroende 1
21565 misstroendeförklaring 1
21566 misstroenderöst 1
21567 misstroendevotum 1
21568 misstrott 1
21569 misstänka 1
21570 misstänker 8
21571 misstänksamhet 3
21572 misstänksamt 1
21573 misstänkt 3
21574 misstänkta 1
21575 misstänkte 3
21576 missuppfattning 2
21577 missuppfattningar 2
21578 missöde 3
21579 missödet 1
21580 mist 3
21581 mista 1
21582 miste 7
21583 mister 1
21584 misär 1
21585 misären 2
21586 mitt 217
21587 mittemot 1
21588 mitten 5
21589 mittgången 1
21590 mittplatsen 1
21591 mix 4
21592 mixas 1
21593 mixtrade 1
21594 mjuk 4
21595 mjuka 3
21596 mjukade 1
21597 mjukare 1
21598 mjukat 1
21599 mjukhjärtad 1
21600 mjuklandning 1
21601 mjukt 1
21602 mjölk 1
21603 mjölke 1
21604 mjölkprodukter 1
21605 mjölkpulver 2
21606 mobilisera 6
21607 mobiliserade 1
21608 mobiliserar 1
21609 mobiliseras 1
21610 mobiliserat 2
21611 mobiliserats 1
21612 mobilisering 3
21613 mobiliseringen 3
21614 mobilområdet 1
21615 mobiltelefoner 2
21616 mobiltelefonerna 1
21617 mobiltelefoni 1
21618 mobiltelefonin 1
21619 mod 8
21620 modebegreppet 1
21621 modell 26
21622 modellen 24
21623 modellens 1
21624 modeller 8
21625 modellerna 4
21626 modenyck 2
21627 modeordet 1
21628 moder 2
21629 moderat 1
21630 moderata 2
21631 modern 11
21632 moderna 21
21633 modernare 1
21634 modernisera 15
21635 moderniserade 1
21636 moderniseras 2
21637 modernisering 38
21638 moderniseringen 5
21639 moderniseringsprocess 2
21640 moderniseringsstrategi 1
21641 modernt 3
21642 moderskap 3
21643 modersmål 1
21644 modet 10
21645 modifiera 1
21646 modifierade 26
21647 modifierat 3
21648 modifierats 1
21649 modig 3
21650 modiga 7
21651 modige 2
21652 modigt 2
21653 modlösa 1
21654 mods 3
21655 modus 2
21656 mogen 3
21657 moget 1
21658 mogna 4
21659 mognad 2
21660 mognat 1
21661 moln 2
21662 molnen 3
21663 molnfria 1
21664 moment 1
21665 momenten 1
21666 momspliktiga 1
21667 monetarism 3
21668 monetaristisk 1
21669 monetaristiska 1
21670 monetär 4
21671 monetära 17
21672 monitoring 1
21673 monokulturer 1
21674 monokulturerna 2
21675 monopol 26
21676 monopolbildning 2
21677 monopolen 1
21678 monopolens 1
21679 monopolet 2
21680 monopolets 1
21681 monopolfrågor 1
21682 monopolföretag 1
21683 monopolföretags 1
21684 monopolintressen 1
21685 monopoliserade 3
21686 monopoliserats 1
21687 monopoliska 1
21688 monopolmarknader 1
21689 monopolrättigheter 1
21690 monopolsituation 1
21691 monopolställning 1
21692 monster 1
21693 monsterhustrun 1
21694 monstermannen 1
21695 monstermasken 1
21696 monsterälskarinnan 1
21697 monterat 1
21698 mor 29
21699 moral 4
21700 moralen 3
21701 moralisk 2
21702 moraliska 7
21703 moraliskt 4
21704 moralism 1
21705 moratorium 1
21706 morbror 17
21707 morbrors 1
21708 mord 10
21709 mordbränder 1
21710 morden 1
21711 mordet 2
21712 mordförsöken 1
21713 mordiska 1
21714 morgnar 1
21715 morgon 120
21716 morgon- 1
21717 morgondagen 2
21718 morgondagens 7
21719 morgonen 4
21720 morgons 1
21721 morgonsolen 1
21722 morgonteet 1
21723 morgontimmen 1
21724 mormodern 1
21725 mormor 3
21726 morot 1
21727 morron 1
21728 morronen 1
21729 mors 2
21730 morse 22
21731 moskiter 1
21732 moskéns 1
21733 moster 6
21734 mot 741
21735 motarbeta 6
21736 motarbetar 1
21737 motbjudande 2
21738 motgångar 1
21739 motgångarna 1
21740 motion 1
21741 motionen 1
21742 motioner 2
21743 motiv 9
21744 motivation 4
21745 motivationen 2
21746 motiven 3
21747 motivera 8
21748 motiverad 2
21749 motiverade 5
21750 motiverades 1
21751 motiverar 9
21752 motiveras 2
21753 motiverat 1
21754 motiverats 1
21755 motivering 7
21756 motiveringar 2
21757 motiveringen 5
21758 motivet 2
21759 motljus 2
21760 motor 3
21761 motorcyklar 3
21762 motorcyklarna 1
21763 motorerna 3
21764 motorindustrin 2
21765 motorister 1
21766 motorn 3
21767 motorns 2
21768 motorväg 2
21769 motorvägar 1
21770 motpart 2
21771 motparten 2
21772 motpartens 1
21773 motparter 1
21774 motpartsmedel 1
21775 motsats 24
21776 motsatsen 11
21777 motsatser 1
21778 motsatsförhållande 1
21779 motsatsställning 1
21780 motsatt 9
21781 motsatta 12
21782 motsatte 2
21783 motstridig 1
21784 motstridiga 8
21785 motstridigheter 2
21786 motsträvig 1
21787 motsträvigt 1
21788 motstycke 6
21789 motstånd 10
21790 motståndare 13
21791 motståndarna 1
21792 motståndet 5
21793 motståndsrörelser 1
21794 motstår 2
21795 motsvara 2
21796 motsvarade 1
21797 motsvarades 1
21798 motsvarande 30
21799 motsvarar 22
21800 motsvaras 1
21801 motsvarats 1
21802 motsvarighet 5
21803 motsvarigheter 2
21804 motsäga 1
21805 motsägande 2
21806 motsägas 1
21807 motsägelse 7
21808 motsägelsefull 1
21809 motsägelsefulla 7
21810 motsägelsefullt 8
21811 motsägelsens 1
21812 motsägelser 3
21813 motsägelserna 1
21814 motsätta 3
21815 motsätter 17
21816 motsättning 8
21817 motsättningar 16
21818 motsättningarna 5
21819 motsättningen 1
21820 motta 1
21821 mottaga 1
21822 mottagande 6
21823 mottagandet 4
21824 mottagare 1
21825 mottagarlandet 2
21826 mottagarlandets 2
21827 mottagarländerna 2
21828 mottagarländernas 1
21829 mottagarna 2
21830 mottagarområden 1
21831 mottagarområdena 1
21832 mottagarprogrammet 1
21833 mottagit 11
21834 mottagits 3
21835 mottagna 1
21836 mottagning 1
21837 mottagningar 1
21838 mottagningsanläggning 1
21839 mottagningsanläggningar 3
21840 mottagningsanläggningen 1
21841 mottagningsanordningar 7
21842 mottagningsanordningarna 1
21843 mottagningsbevis 1
21844 mottagningsceremoni 1
21845 mottagningsförhållanden 1
21846 mottar 1
21847 motto 1
21848 mottog 3
21849 mottogs 1
21850 motverka 9
21851 motverkar 2
21852 motvikt 2
21853 motvilligt 3
21854 motvärn 1
21855 motåtgärd 1
21856 motåtgärder 5
21857 moçambikier 2
21858 moçambikierna 1
21859 moçambikiska 3
21860 mr 22
21861 mrs 13
21862 muddermassorna 1
21863 muddras 1
21864 mugglare 2
21865 mugglarkvinna 1
21866 mugglarpengar 1
21867 mugglarägare 1
21868 mullrande 1
21869 multi-etniska 1
21870 multi-etniskt 1
21871 multietnisk 1
21872 multietniska 3
21873 multietniskt 2
21874 multilateral 2
21875 multilaterala 7
21876 multinationell 1
21877 multinationella 15
21878 multinationellt 1
21879 multipliceras 1
21880 multiplikatoreffekt 2
21881 multiplikatoreffekten 1
21882 mumifierade 1
21883 mumla 1
21884 mumlade 3
21885 mumlande 1
21886 mun 4
21887 munnen 5
21888 munterhet 1
21889 muntert 1
21890 muntlig 2
21891 muntliga 23
21892 muntligen 1
21893 muntligt 4
21894 muntra 1
21895 mur 2
21896 murad 1
21897 murar 3
21898 museifartyg 1
21899 museifartygen 1
21900 muselmansk 1
21901 museum 1
21902 musik 5
21903 musikanter 1
21904 musiken 3
21905 musiker 1
21906 muskler 1
21907 muskulös 1
21908 muslim 1
21909 mussel- 3
21910 musselodlare 2
21911 must 1
21912 mustasch 1
21913 mustascherna 1
21914 muta 1
21915 mutor 1
21916 muttrade 3
21917 muttrande 2
21918 mycken 3
21919 mycket 1390
21920 mygg 1
21921 myggen 1
21922 myggor 1
21923 myllan 1
21924 myllrade 2
21925 myllrande 1
21926 myllrar 1
21927 myndiga 1
21928 myndigförklarade 1
21929 myndighet 27
21930 myndigheten 30
21931 myndighetens 16
21932 myndigheter 68
21933 myndigheterna 105
21934 myndigheternas 13
21935 myndigheters 4
21936 myndighetsförfaranden 1
21937 myndighetskrångel 1
21938 myndighetsåtgärder 1
21939 mynna 4
21940 mynning 2
21941 mynningarna 1
21942 mynningen 3
21943 mynningsområde 1
21944 mynningsområdet 1
21945 mynt 4
21946 mynten 2
21947 myror 2
21948 mysteriejakt 1
21949 mysterier 1
21950 mysterium 4
21951 mystiska 2
21952 mytiskt 1
21953 mäkleriverksamhet 1
21954 mäkta 1
21955 mäktig 1
21956 mäktiga 2
21957 mäktigaste 1
21958 män 76
21959 mängd 33
21960 mängden 7
21961 mängder 11
21962 mängdfunktionerna 1
21963 mängdfunktionsreferens 1
21964 männen 20
21965 männens 3
21966 människa 14
21967 människan 14
21968 människans 9
21969 människo- 1
21970 människoben 1
21971 människoföda 2
21972 människoföraktande 1
21973 människoförföljande 1
21974 människohandel 3
21975 människoknotor 1
21976 människokompost 1
21977 människokännedom 1
21978 människokärlek 1
21979 människoliv 10
21980 människomassan 1
21981 människomyller 1
21982 människonaglar 1
21983 människor 213
21984 människorna 50
21985 människornas 5
21986 människors 35
21987 människorätten 1
21988 människorättskommissionerna 1
21989 människorättsnarcissismen 1
21990 människorättsnivån 1
21991 människorättsorganisationer 2
21992 människorättspolitik 5
21993 människorättspolitiken 3
21994 människosläktet 2
21995 människosmugglarnas 1
21996 människosmuggling 1
21997 människosyn 1
21998 människovänlig 1
21999 människovärdet 1
22000 människovärdiga 2
22001 människovärdigt 1
22002 mäns 2
22003 mänsklig 15
22004 mänskliga 247
22005 mänskligheten 6
22006 mänskligt 6
22007 märk 1
22008 märka 6
22009 märkas 1
22010 märkbar 5
22011 märkbara 3
22012 märkbart 2
22013 märke 16
22014 märken 5
22015 märker 4
22016 märkesgrupperna 1
22017 märklig 3
22018 märkliga 3
22019 märkligare 1
22020 märkligheter 1
22021 märkligt 4
22022 märkning 13
22023 märkningen 4
22024 märks 1
22025 märkt 2
22026 märkte 3
22027 märkvärdig 1
22028 märkvärdiga 1
22029 märkvärdigt 4
22030 mäss 1
22031 mässingsinstrument 1
22032 mästerverk 2
22033 mäta 7
22034 mätare 3
22035 mätas 5
22036 mätbara 2
22037 mäter 1
22038 mätningar 1
22039 mäts 3
22040 mätt 2
22041 mätte 1
22042 må 17
22043 måfå 1
22044 måhända 7
22045 mål 282
22046 mål-2-området 1
22047 måla 3
22048 målade 3
22049 målar 1
22050 målarfärg 1
22051 målas 1
22052 målat 1
22053 målats 2
22054 målen 47
22055 målens 1
22056 målet 62
22057 målformat 1
22058 målgrupp 2
22059 målgrupper 1
22060 målgången 1
22061 målinriktad 1
22062 målinriktade 2
22063 målinriktat 5
22064 mållösa 1
22065 målmedvetet 3
22066 målområdena 1
22067 målområdet 1
22068 målsättning 25
22069 målsättningar 25
22070 målsättningarna 16
22071 målsättningen 16
22072 måltid 2
22073 måltidens 1
22074 mån 31
22075 mån. 1
22076 måna 3
22077 månad 33
22078 månaden 16
22079 månader 89
22080 månaderna 34
22081 månaders 1
22082 månads 2
22083 månadslånga 1
22084 månadsvisa 1
22085 månatliga 1
22086 månbelyst 1
22087 måndag 7
22088 måndagar 1
22089 måndagen 2
22090 måndags 11
22091 månde 1
22092 måne 1
22093 många 559
22094 mångbesjungna 1
22095 mångfald 25
22096 mångfalden 16
22097 mångfaldig 1
22098 mångfaldiga 4
22099 mångfaldigandet 1
22100 mångfaldigas 1
22101 mångfaldigt 2
22102 mångformiga 1
22103 mångfunktionell 1
22104 mångfärgad 1
22105 mångkulturella 2
22106 mångkunnig 1
22107 mångnationellt 1
22108 mångsidighet 1
22109 mångsidigt 4
22110 mångskiftande 1
22111 mångt 2
22112 mångtaliga 1
22113 mångtydiga 1
22114 mångåriga 2
22115 månljuset 1
22116 månsken 1
22117 mår 3
22118 måste 1948
22119 mått 9
22120 måtte 2
22121 måttenhet 1
22122 måttet 1
22123 måttfulla 1
22124 måttfullhet 1
22125 måttlig 1
22126 måtto 7
22127 måttstock 4
22128 måttstocken 1
22129 möblemanget 1
22130 möbler 3
22131 möblerad 1
22132 möblerna 1
22133 möda 5
22134 mödan 1
22135 mödosam 1
22136 mödosamma 1
22137 mödosamt 1
22138 mödrar 2
22139 möjlig 15
22140 möjliga 63
22141 möjligen 12
22142 möjliggjorde 1
22143 möjliggjort 3
22144 möjliggör 13
22145 möjliggöra 23
22146 möjliggörs 2
22147 möjlighet 130
22148 möjligheten 54
22149 möjligheter 129
22150 möjligheterna 22
22151 möjligheternas 4
22152 möjligheteten 1
22153 möjligt 335
22154 möjligtvis 3
22155 mönster 4
22156 mönsterbild 1
22157 mönsterskydd 1
22158 mönstring 1
22159 mördade 1
22160 mördades 2
22161 mördande 2
22162 mördar 1
22163 mördare 1
22164 mördaren 1
22165 mördas 1
22166 mördat 2
22167 mördats 2
22168 mörk 4
22169 mörka 16
22170 mörkare 2
22171 mörkblond 1
22172 mörkblå 1
22173 mörker 4
22174 mörklägga 1
22175 mörknade 1
22176 mörkret 12
22177 mörkrets 1
22178 mörkrött 1
22179 mörkt 6
22180 möta 26
22181 möte 46
22182 möten 14
22183 mötena 2
22184 möter 7
22185 mötes 6
22186 mötespunkt 1
22187 mötet 22
22188 möts 3
22189 mött 1
22190 mötte 1
22191 möttes 3
22192 mötts 1
22193 müssen 2
22194 n 2
22195 nackdel 8
22196 nackdelar 7
22197 nacken 4
22198 nagel 1
22199 naglar 1
22200 naiva 1
22201 naivitet 1
22202 naivt 1
22203 nakna 2
22204 nallebjörn 1
22205 namn 49
22206 namnen 1
22207 namnet 23
22208 namnfrågan 1
22209 namnlös 1
22210 namnlösa 1
22211 namnteckning 2
22212 namnupprop 6
22213 nappat 1
22214 narkotika 3
22215 narkotikabekämpning 1
22216 narkotikahandel 1
22217 narkotikahandeln 1
22218 narkotikamissbrukare 1
22219 narkotikan 1
22220 narkotikaproblematiken 1
22221 narkotikasmuggling 2
22222 narrarnas 1
22223 nation 5
22224 national 1
22225 national-socialistiska 1
22226 nationalekonomin 1
22227 nationalekonomisk 1
22228 nationalekonomiska 3
22229 nationalekonomiskt 2
22230 nationalförsamling 1
22231 nationalförsamlingen 3
22232 nationaliseringsprocess 1
22233 nationalism 4
22234 nationalismens 1
22235 nationalister 1
22236 nationalisterna 1
22237 nationalistiska 1
22238 nationalitet 5
22239 nationaliteter 3
22240 nationalliberaler 1
22241 nationalräkenskapssystemet 6
22242 nationalsocialismen 1
22243 nationalstaten 2
22244 nationalstatens 1
22245 nationalstater 2
22246 nationalstaterna 1
22247 nationell 46
22248 nationella 260
22249 nationellt 13
22250 nationen 1
22251 nationens 2
22252 nationer 12
22253 nationerna 25
22254 nationernas 39
22255 nationsgränser 2
22256 nationsregionerna 1
22257 nationsskapande 1
22258 nationsspecifika 1
22259 natt 3
22260 nattblommor 1
22261 natten 15
22262 nattens 1
22263 nattetid 1
22264 nattfjärilar 1
22265 nattfjärilsmjuka 1
22266 nattliga 2
22267 nattlinne 1
22268 nattsammanträden 1
22269 nattsammanträdenas 1
22270 nattsäck 1
22271 nattupplagan 1
22272 nattvagabonderande 1
22273 nattvinden 1
22274 nattväskan 1
22275 natur 29
22276 natur- 3
22277 natura 1
22278 naturarvet 1
22279 naturen 18
22280 naturens 2
22281 naturfenomen 1
22282 naturkatastrof 2
22283 naturkatastrofen 2
22284 naturkatastrofer 17
22285 naturlig 7
22286 naturliga 19
22287 naturligt 16
22288 naturligtvis 237
22289 naturnätverket 1
22290 naturnödvändighet 1
22291 naturområden 2
22292 naturresurs 3
22293 naturresurser 4
22294 naturresurserna 5
22295 naturskydd 1
22296 naturskyddspolitiken 1
22297 naturtillgångar 4
22298 naturvetenskaplig 1
22299 naturvidrigt 1
22300 navajoindianerna 1
22301 navajoreservatet 1
22302 navigationssektionen 1
22303 navigerat 1
22304 nazism 2
22305 nazismen 4
22306 nazismens 1
22307 nazist 2
22308 nazistflirtande 1
22309 nazistisk 1
22310 ne 1
22311 necessär 2
22312 necessären 1
22313 ned 65
22314 nedan 1
22315 nedanför 4
22316 nedbrytningen 1
22317 nedbrända 1
22318 nedbäddad 1
22319 neddragna 1
22320 neddragningar 1
22321 nederbörd 1
22322 nederbörden 2
22323 nederlag 2
22324 nederländare 1
22325 nederländsk 11
22326 nederländsk-brittisk-skandinavisk 1
22327 nederländska 15
22328 nedersta 1
22329 nedför 1
22330 nedgång 3
22331 nedgången 2
22332 nedifrån 1
22333 nedkomma 1
22334 nedkomst 1
22335 nedlagd 1
22336 nedlagda 1
22337 nedläggning 2
22338 nedläggningar 2
22339 nedläggningen 1
22340 nedlåta 1
22341 nedlåtande 1
22342 nedmontera 1
22343 nedmontering 2
22344 nedmonterings- 1
22345 nedrullningsbara 1
22346 nedrustning 1
22347 nedrustningen 1
22348 nedskräpningsproblem 1
22349 nedskärning 2
22350 nedskärningar 6
22351 nedskärningspolitik 1
22352 nedsmutsade 2
22353 nedsmutsning 3
22354 nedsmutsningen 4
22355 nedströms 5
22356 nedstämd 1
22357 nedstängning 1
22358 nedstängningsplaner 1
22359 nedsättande 1
22360 nedtecknat 1
22361 nedvärdera 1
22362 nedvärderas 1
22363 nedåt 6
22364 negativ 14
22365 negativa 38
22366 negativism 1
22367 negativt 21
22368 neger 1
22369 negligera 1
22370 nej 25
22371 nejlikor 1
22372 neka 3
22373 nekad 1
22374 nekande 1
22375 nekas 5
22376 neo-liberalism 1
22377 neofascistiska 2
22378 neoklassiska 1
22379 neokolonial 1
22380 neokolonialismen 1
22381 neokolonialistiska 1
22382 neonazistiskt 1
22383 neonlampor 1
22384 nepotism 5
22385 ner 81
22386 nerdrogad 1
22387 nere 16
22388 nerför 9
22389 nerhukade 1
22390 nerver 1
22391 nervkrig 1
22392 nervpåfrestande 1
22393 nervös 2
22394 nervösa 1
22395 nervöst 1
22396 nettoupplåning 1
22397 nettoökning 1
22398 neutral 1
22399 neutrala 2
22400 neutraliserar 1
22401 neutraliseras 1
22402 neutralitet 1
22403 neutralt 2
22404 neutre 2
22405 new 6
22406 ni 825
22407 nickade 1
22408 nigerianska 1
22409 nihilo-rätt 1
22410 nikotinproblemen 1
22411 nimbus 1
22412 nio 17
22413 nionde 2
22414 nioåring 1
22415 nischer 1
22416 nit 1
22417 nitratdirektivet 1
22418 nittiotalet 1
22419 nitton 2
22420 nittonhundra 1
22421 nittonhundrafyrtitalet 1
22422 nittonhundratalet 1
22423 nittonhundratalets 1
22424 nivå 168
22425 nivåer 23
22426 nivåerna 2
22427 nivån 15
22428 njuta 2
22429 njuter 2
22430 njutning 1
22431 njöt 3
22432 nn 1
22433 no 6
22434 nobelpristagaren 1
22435 nog 53
22436 noga 35
22437 noggrann 7
22438 noggranna 5
22439 noggrannare 4
22440 noggrannhet 4
22441 noggrannheten 1
22442 noggrant 28
22443 noll 17
22444 noll-alternativet 1
22445 nollgradig 3
22446 nollgränsvärde 1
22447 nollkravet 1
22448 nollning 1
22449 nollnivå 1
22450 nollnivårisk 1
22451 nollor 1
22452 nollrisk 1
22453 nollstrecket 1
22454 nollställda 1
22455 nollutsläpp 2
22456 nollårig 1
22457 nominell 2
22458 nominella 2
22459 nominera 4
22460 nominerade 1
22461 nominerar 1
22462 nomineras 1
22463 nomineringen 1
22464 non 4
22465 nonchalansen 1
22466 nonchalant 1
22467 nonchalerade 2
22468 nonsens 1
22469 nonsensord 1
22470 nord 1
22471 nord-syd 2
22472 nordafrikanska 3
22473 nordamerikanerna 1
22474 nordamerikanska 6
22475 nordeuropeiska 1
22476 nordirländare 1
22477 nordirländska 1
22478 nordisk 1
22479 nordiska 4
22480 nordkusten 1
22481 nordlig 1
22482 nordliga 6
22483 nordtyska 1
22484 nordvästra 4
22485 norm 2
22486 normal 5
22487 normala 9
22488 normaliserades 1
22489 normalisering 5
22490 normaliseringen 2
22491 normalitet 1
22492 normalt 17
22493 normativ 1
22494 normativt 2
22495 normen 1
22496 normer 36
22497 normerna 15
22498 normgivande 1
22499 norr 9
22500 norr-söder 1
22501 norra 25
22502 norrmännens 1
22503 norrut 2
22504 norska 2
22505 norskt 1
22506 nos 1
22507 noshörning 1
22508 nostrum 1
22509 not 2
22510 notan 1
22511 notera 23
22512 noterade 6
22513 noterades 1
22514 noterar 28
22515 noteras 3
22516 noterat 17
22517 noterna 1
22518 notis 1
22519 november 30
22520 nr 81
22521 nu 697
22522 nuet 1
22523 nuets 1
22524 null-värden 5
22525 nulla 1
22526 nullitetssanktionen 1
22527 nullvärde 1
22528 nuläget 5
22529 numer 1
22530 numera 19
22531 numerära 1
22532 nummer 11
22533 numreringen 1
22534 numret 6
22535 nunnor 1
22536 nutida 1
22537 nuvarande 141
22538 ny 173
22539 nya 621
22540 nyanlända 1
22541 nyansera 1
22542 nyanserad 1
22543 nyanserna 1
22544 nyanställda 2
22545 nyanställningar 1
22546 nyare 1
22547 nyaste 1
22548 nybildande 1
22549 nybilsköparna 1
22550 nybilspriset 1
22551 nybyggets 1
22552 nyckel 1
22553 nyckelfaktor 1
22554 nyckelfråga 3
22555 nyckelfrågan 1
22556 nyckelfrågor 1
22557 nyckelfrågorna 1
22558 nyckelfunktioners 1
22559 nyckeln 6
22560 nyckelområden 1
22561 nyckelord 1
22562 nyckelorden 1
22563 nyckelordet 1
22564 nyckelproblem 2
22565 nyckelpunkter 1
22566 nyckelroll 3
22567 nyckelsektor 1
22568 nyckelåtgärder 1
22569 nycklar 1
22570 nycklarna 1
22571 nydanande 6
22572 nye 3
22573 nyetableringar 1
22574 nyexaminerad 1
22575 nyfascister 1
22576 nyfattigdom 1
22577 nyfiken 4
22578 nyfiket 1
22579 nyfikna 1
22580 nyföretagarvänlig 1
22581 nyförvärvade 1
22582 nygift 1
22583 nyhet 6
22584 nyheten 1
22585 nyheter 14
22586 nyheterna 9
22587 nyhetsinslag 1
22588 nyhetsprogrammet 1
22589 nyhetsrapporterna 1
22590 nykomlingar 1
22591 nykomlingarna 1
22592 nyktert 3
22593 nyktra 1
22594 nylansera 1
22595 nylansering 1
22596 nylanseringen 1
22597 nyliberal 2
22598 nyliberala 2
22599 nyliberalt 1
22600 nyligen 84
22601 nylon 1
22602 nylonet 1
22603 nylonspetsar 1
22604 nylontrosornas 1
22605 nynazism 1
22606 nynazismen 1
22607 nynazist 1
22608 nynazister 2
22609 nynazistiska 1
22610 nypa 1
22611 nypan 1
22612 nyplanteringen 1
22613 nyskapande 3
22614 nyss 46
22615 nystart 1
22616 nytt 152
22617 nytta 53
22618 nyttan 5
22619 nyttig 7
22620 nyttiga 8
22621 nyttighet 1
22622 nyttigt 4
22623 nyttjande 1
22624 nyttoanalys 1
22625 nyttobruk 1
22626 nyttofordon 9
22627 nytänkande 3
22628 nyval 1
22629 nyvald 1
22630 nyvalda 1
22631 nyvalde 1
22632 nyårsaftonen 1
22633 nämligen 204
22634 nämna 63
22635 nämnare 1
22636 nämnaren 2
22637 nämnas 3
22638 nämnda 16
22639 nämnde 45
22640 nämndes 9
22641 nämner 24
22642 nämns 23
22643 nämnt 26
22644 nämnts 20
22645 nämnvärd 1
22646 nämnvärda 1
22647 nämnvärt 1
22648 när 1068
22649 nära 79
22650 närapå 1
22651 närbelägna 2
22652 närbesläktad 1
22653 närbesläktade 1
22654 närekonomi 1
22655 närhelst 1
22656 närhet 1
22657 närheten 14
22658 närhetsamtal 1
22659 näring 1
22660 näringar 3
22661 näringsgren 3
22662 näringsgrenen 1
22663 näringsidkare 1
22664 näringskedja 1
22665 näringskedjan 1
22666 näringsliv 1
22667 näringslivet 14
22668 näringslivets 5
22669 näringslivsaktörer 1
22670 näringsrik 1
22671 näringsstrukturen 1
22672 näringstillskott 1
22673 näringsvärden 1
22674 närliggande 1
22675 närma 10
22676 närmade 2
22677 närmande 10
22678 närmanden 1
22679 närmandet 1
22680 närmar 8
22681 närmare 50
22682 närmast 16
22683 närmaste 53
22684 närmsta 1
22685 närområdet 2
22686 närpolisen 1
22687 närpoliser 1
22688 närpolissystem 1
22689 närstående 4
22690 närsynt 2
22691 närvara 6
22692 närvarade 1
22693 närvarande 123
22694 närvarar 1
22695 närvaro 25
22696 närvaron 5
22697 näsa 4
22698 näsan 8
22699 näsborrar 1
22700 näsdukar 1
22701 näsduken 1
22702 näst 1
22703 nästa 96
22704 nästan 86
22705 nästkommande 1
22706 näsvingarna 1
22707 nät 12
22708 näten 5
22709 nätens 1
22710 nätet 3
22711 nätstrukturer 1
22712 nätt 2
22713 nätter 2
22714 nätterna 1
22715 nätverk 13
22716 nätverken 3
22717 nätverkens 2
22718 nätverket 2
22719 nätverkslicens 1
22720 nätverkslicensavtal 1
22721 nätverkslicensen 1
22722 nätverkssamhället 1
22723 nå 70
22724 nåbar 2
22725 nåd 2
22726 nådde 5
22727 nåddes 2
22728 nåden 1
22729 någon 445
22730 någons 1
22731 någonsin 30
22732 någonstans 24
22733 någonting 108
22734 någonvart 1
22735 någorlunda 2
22736 något 612
22737 någotdera 1
22738 några 453
22739 nåja 1
22740 nål 1
22741 nån 3
22742 nånsin 3
22743 nånstans 4
22744 nånting 3
22745 når 9
22746 nås 4
22747 nåt 5
22748 nått 21
22749 nåtts 1
22750 nöd 3
22751 nödbedd 1
22752 nöden 2
22753 nödens 1
22754 nödfall 1
22755 nödgas 2
22756 nödhjälp 4
22757 nödhjälpen 1
22758 nödinsatser 1
22759 nödlösning 1
22760 nödraketer 1
22761 nödreparationer 1
22762 nödsituation 2
22763 nödsituationen 1
22764 nödsituationer 1
22765 nödsituationsfasen 1
22766 nödställda 1
22767 nödtorftiga 1
22768 nödvändig 51
22769 nödvändiga 85
22770 nödvändigare 1
22771 nödvändiggör 1
22772 nödvändighet 12
22773 nödvändigheten 18
22774 nödvändigheterna 1
22775 nödvändighetsperspektiv 1
22776 nödvändigt 205
22777 nödvändigtvis 18
22778 nödåtgärder 1
22779 nöja 20
22780 nöjaktig 1
22781 nöjaktigt 1
22782 nöjd 14
22783 nöjda 16
22784 nöjde 1
22785 nöje 12
22786 nöjer 6
22787 nöjesbåtar 1
22788 nöjet 6
22789 nöjsam 1
22790 nöjt 2
22791 nöt 1
22792 nötkreatur 1
22793 nötkött 6
22794 nötkötts- 1
22795 nötköttsöverskott 1
22796 nötskal 2
22797 nött 1
22798 nötter 1
22799 nötterna 1
22800 nöttköttslager 1
22801 o 3
22802 o.s.v. 2
22803 oacceptabel 18
22804 oacceptabelt 30
22805 oacceptabla 17
22806 oaktat 2
22807 oanmälda 3
22808 oansenligt 1
22809 oanständiga 1
22810 oansvariga 3
22811 oansvarighet 6
22812 oansvarigheten 1
22813 oanvända 1
22814 oanvändbar 2
22815 oanvändbart 1
22816 oartig 1
22817 oavbruten 2
22818 oavbrutet 2
22819 oavbrutna 1
22820 oavhängighet 2
22821 oavhängighetsförklaringen 2
22822 oavsett 41
22823 oavsiktlig 1
22824 oavsiktliga 3
22825 oavsiktligt 1
22826 oavslutade 1
22827 oavvislig 1
22828 obalans 6
22829 obalansen 5
22830 obalanser 2
22831 obalanserna 2
22832 obarmhärtiga 1
22833 obarmhärtigt 1
22834 obeboelig 1
22835 obefintliga 2
22836 obefläckad 2
22837 obefogat 2
22838 obegriplig 2
22839 obegripliga 1
22840 obegripligt 3
22841 obegränsad 6
22842 obegränsat 1
22843 obehag 1
22844 obehagliga 2
22845 obehagligt 4
22846 obekant 1
22847 obekanta 1
22848 obekväma 1
22849 obekymrade 1
22850 obemannad 1
22851 obemärkt 2
22852 obemärkthet 1
22853 oberoende 83
22854 oberoendes 1
22855 oberoendet 1
22856 oberättigad 1
22857 oberättigat 1
22858 oberörd 2
22859 oberörda 1
22860 obestridlig 1
22861 obestridliga 2
22862 obestämd 4
22863 obesvarad 1
22864 obesvarade 3
22865 obesvärade 1
22866 obetalda 2
22867 obetydlig 2
22868 obetydligt 1
22869 obevakade 1
22870 obevekliga 1
22871 obeveklighet 1
22872 obeväpnade 1
22873 obildad 1
22874 objekt 5
22875 objektbibliotek 1
22876 objektdefinitioner 1
22877 objektet 2
22878 objektets 1
22879 objektiv 3
22880 objektiva 5
22881 objektivt 7
22882 oblandad 1
22883 obligationer 1
22884 obligationsmarknaderna 1
22885 obligatorisk 13
22886 obligatoriska 12
22887 obligatoriskt 4
22888 obligatorium 1
22889 obrukbart 1
22890 observation 1
22891 observationerna 1
22892 observatorium 1
22893 observatory 2
22894 observatörens 1
22895 observatörer 6
22896 observatörerna 1
22897 observera 2
22898 observerats 1
22899 obsolet 1
22900 obundna 3
22901 oceanen 1
22902 oceanerna 2
22903 oceanernas 1
22904 och 15193
22905 också 1574
22906 ockupanten 1
22907 ockupation 2
22908 ockupationen 4
22909 ockupationsmakt 1
22910 ockupationsstyrkorna 1
22911 ockuperade 15
22912 ockuperades 1
22913 ockuperande 1
22914 ockuperas 1
22915 ockuperat 1
22916 odds 1
22917 odefinierade 1
22918 odefinierbart 1
22919 odelad 1
22920 odelade 1
22921 odelbara 1
22922 odemokratiska 2
22923 odiskutabel 1
22924 odiskutabelt 1
22925 odjur 2
22926 odla 4
22927 odlad 1
22928 odlar 1
22929 odlare 1
22930 odlarna 3
22931 odling 3
22932 odlingar 7
22933 odlingarna 1
22934 odlingen 1
22935 odlingsmarker 1
22936 odlingsplatser 1
22937 odugliga 1
22938 odödliga 1
22939 oeftergivligt 1
22940 oegennyttiga 2
22941 oegentlig 1
22942 oegentliga 1
22943 oegentlighet 2
22944 oegentligheter 3
22945 oegentligheterna 1
22946 oegentligt 1
22947 oekonomisk 1
22948 oekonomiskt 1
22949 oemotståndlig 1
22950 oemotståndligt 1
22951 oemotsägligt 1
22952 oenighet 5
22953 oenigheten 1
22954 oenigheterna 1
22955 oense 5
22956 oerhörd 4
22957 oerhörda 5
22958 oerhört 25
22959 oersättliga 1
22960 oetiska 1
22961 of 11
22962 ofantlig 1
22963 ofantliga 5
22964 ofantligt 1
22965 ofarlig 2
22966 ofarligt 1
22967 ofattbara 3
22968 ofattbart 1
22969 ofelbara 1
22970 offensiv 2
22971 offensiva 1
22972 offensiven 1
22973 offensivt 3
22974 offentlig 38
22975 offentliga 152
22976 offentligen 1
22977 offentliggjorda 1
22978 offentliggjorde 5
22979 offentliggjordes 2
22980 offentliggjort 3
22981 offentliggjorts 4
22982 offentliggör 2
22983 offentliggöra 7
22984 offentliggörande 1
22985 offentliggörandet 2
22986 offentliggöras 6
22987 offentliggörs 5
22988 offentlighet 2
22989 offentligheten 2
22990 offentlighetens 2
22991 offentlighetsförordningen 1
22992 offentlighetskampanj 1
22993 offentlighetsprincip 1
22994 offentligpolitiska 1
22995 offentligt 16
22996 offer 32
22997 officerare 1
22998 officiell 1
22999 officiella 18
23000 officiellt 5
23001 offra 1
23002 offrade 1
23003 offrades 1
23004 offrar 1
23005 offras 4
23006 offren 25
23007 offrens 4
23008 offret 2
23009 oflexibilitet 1
23010 oformaterad 1
23011 oframkomlig 1
23012 ofred 1
23013 ofruktbart 1
23014 ofrånkomligen 3
23015 ofrånkomligt 3
23016 ofta 157
23017 oftare 14
23018 oftast 7
23019 ofullkomlighet 1
23020 ofullkomligt 1
23021 ofullständig 3
23022 ofullständiga 4
23023 ofullständigt 1
23024 ofärdig 1
23025 oförblommerat 1
23026 ofördelaktiga 1
23027 ofördelaktigaste 1
23028 ofördelaktigt 2
23029 oförenlig 2
23030 oförenliga 2
23031 oförenlighet 1
23032 oförenligt 4
23033 oförklarat 1
23034 oförklarlig 2
23035 oförklarligt 1
23036 oförlåtlig 1
23037 oförlåtligt 1
23038 oförmåga 7
23039 oförmågan 3
23040 oförmögen 3
23041 oförmögna 1
23042 oförnekligen 1
23043 oförnuftigt 1
23044 oförorenade 1
23045 oförsiktigt 1
23046 oförskämda 1
23047 oförståeligt 2
23048 oförsvarlig 2
23049 oförsvarligt 1
23050 oförtjänt 1
23051 oförtrutet 1
23052 oförtröttat 1
23053 oförutsägbar 1
23054 oföränderlig 2
23055 oföränderliga 1
23056 oföränderlighet 1
23057 oförändrad 2
23058 oförändrade 4
23059 oförändrat 1
23060 ogenomförbar 2
23061 ogenomskinligheten 1
23062 ogenomträngligt 1
23063 ogifta 1
23064 ogillande 1
23065 ogrundad 1
23066 ogrundat 1
23067 ogräs 1
23068 ogynnsam 1
23069 ogynnsamma 2
23070 ogynnsamt 1
23071 ohejdad 1
23072 ohjälpligt 2
23073 ohyggliga 1
23074 ohyggligt 1
23075 ohygienisk 2
23076 ohyra 1
23077 ohälsa 1
23078 ohälsosamma 2
23079 ohälsosamt 1
23080 ohämmad 2
23081 ohämmade 3
23082 ohållbar 1
23083 ohållbara 1
23084 ohållbart 1
23085 ohörsamma 1
23086 ohövlig 2
23087 ohövliga 1
23088 oigenkännelighet 1
23089 oinskränkt 1
23090 oinskränkta 2
23091 oinspelade 1
23092 ointelligent 1
23093 ointressant 1
23094 ointresse 3
23095 ointresserad 1
23096 ointresset 1
23097 ojämförbar 1
23098 ojämlik 1
23099 ojämlikhet 9
23100 ojämlikheten 3
23101 ojämlikheter 3
23102 ojämlikheterna 1
23103 ojämn 1
23104 ojämna 2
23105 ojämnt 3
23106 okaraktäristiskt 1
23107 oket 1
23108 oklanderlig 2
23109 oklanderliga 1
23110 oklanderligt 1
23111 oklar 4
23112 oklara 4
23113 oklarhet 4
23114 oklarheter 5
23115 oklart 5
23116 oklok 1
23117 oklokt 1
23118 okomplicerad 1
23119 okomplicerade 2
23120 okonstlad 1
23121 okontrollerad 4
23122 okontrollerade 3
23123 okontrollerat 1
23124 okontrollerbar 1
23125 okontrollerbara 1
23126 okritiska 1
23127 okritiskt 3
23128 okränkbara 2
23129 okränkbarheten 1
23130 oktaverna 1
23131 oktober 24
23132 okunnig 3
23133 okunniga 1
23134 okunnighet 6
23135 okunnigt 1
23136 okunskap 1
23137 okuvlig 1
23138 okänd 1
23139 okända 4
23140 okänslig 1
23141 okänsliga 1
23142 okänt 1
23143 olaglig 1
23144 olagliga 3
23145 olagligheter 2
23146 olagligt 5
23147 olet 1
23148 olidliga 1
23149 oligarki 1
23150 oligarkier 1
23151 olik 1
23152 olika 436
23153 olikartade 2
23154 olikhet 1
23155 olikheter 8
23156 olikheterna 4
23157 oliver 2
23158 olja 11
23159 oljan 7
23160 oljebefraktaren 1
23161 oljeblanka 2
23162 oljebolag 2
23163 oljebolagen 4
23164 oljebolagens 2
23165 oljebolaget 2
23166 oljebälte 7
23167 oljebälten 2
23168 oljebältena 1
23169 oljebältet 7
23170 oljebältets 1
23171 oljeeldningen 1
23172 oljefartyg 4
23173 oljefartygen 1
23174 oljefläckar 1
23175 oljeföroreningar 2
23176 oljeföroreningarna 2
23177 oljeföroreningens 1
23178 oljeindränkta 3
23179 oljeindustrin 1
23180 oljeinkomsterna 1
23181 oljekoka 1
23182 oljekoncernerna 1
23183 oljekontrakt 1
23184 oljelast 1
23185 oljepriser 1
23186 oljeproducenterna 1
23187 oljerester 1
23188 oljeskadefonderna 1
23189 oljeslam 2
23190 oljespill 1
23191 oljestället 1
23192 oljetankbåtar 1
23193 oljetankern 3
23194 oljetankerns 2
23195 oljetankfartyg 2
23196 oljetankfartyget 1
23197 oljetankrar 2
23198 oljetankrarna 1
23199 oljetankrarnas 1
23200 oljetransporter 1
23201 oljetrusterna 1
23202 oljeutsläpp 5
23203 oljeutsläppen 1
23204 oljeutsläppet 1
23205 oljeutvinningsplattformar 1
23206 oljevägen 1
23207 oljig 1
23208 oljiga 2
23209 ologiska 1
23210 olycka 19
23211 olyckan 7
23212 olycklig 5
23213 olyckliga 9
23214 olyckligt 4
23215 olyckligtvis 1
23216 olyckor 20
23217 olyckorna 1
23218 olycksbringande 1
23219 olycksbådande 2
23220 olycksdiger 1
23221 olycksdrabbade 5
23222 olycksfall 1
23223 olycksfallsförsäkringar 1
23224 olycksfåglar 1
23225 olyckshändelse 1
23226 olyckshändelsen 1
23227 olycksrisker 1
23228 olycksriskerna 1
23229 olycksöde 1
23230 olydig 1
23231 olympiska 1
23232 olägenhetslagstiftningarna 1
23233 olämplig 2
23234 olämpliga 3
23235 olämpligt 5
23236 olösligt 1
23237 olösta 3
23238 om 5768
23239 omarbetning 2
23240 ombads 3
23241 ombeds 2
23242 ombesörja 4
23243 ombesörjer 1
23244 ombetts 2
23245 ombonat 1
23246 ombord 9
23247 ombud 2
23248 ombuden 1
23249 ombudsmannen 7
23250 ombudsmannens 8
23251 ombyggnad 1
23252 ombytligt 1
23253 omcentrera 1
23254 omdebatterade 1
23255 omdefiniera 2
23256 omdefinieras 1
23257 omdefiniering 1
23258 omdirigerade 1
23259 omdirigerades 1
23260 omdirigerar 1
23261 omdirigeras 1
23262 omdirigering 1
23263 omdiskuterade 1
23264 omdöme 3
23265 omdömesförmåga 2
23266 omdömesgilla 1
23267 omedelbar 7
23268 omedelbara 5
23269 omedelbart 44
23270 omedgörlig 2
23271 omedveten 1
23272 omedvetet 3
23273 omen 1
23274 omfatta 42
23275 omfattade 1
23276 omfattades 3
23277 omfattande 87
23278 omfattar 53
23279 omfattas 33
23280 omfattning 20
23281 omfattningen 8
23282 omflyttning 2
23283 omflyttningar 2
23284 omflyttningen 1
23285 omforma 1
23286 omformulerad 1
23287 omformulerar 1
23288 omformuleras 1
23289 omformulering 2
23290 omfånget 2
23291 omfångsrikt 1
23292 omfördelande 1
23293 omfördelning 5
23294 omfördelningen 2
23295 omförhandlingen 1
23296 omge 1
23297 omger 3
23298 omges 2
23299 omgestaltandet 1
23300 omgift 1
23301 omgivande 3
23302 omgiven 1
23303 omgivet 1
23304 omgivna 1
23305 omgivning 3
23306 omgivningar 1
23307 omgivningarna 1
23308 omgivningen 2
23309 omgruppera 1
23310 omgrupperingar 1
23311 omgående 2
23312 omgång 2
23313 omgångarna 1
23314 omgången 5
23315 omhulda 1
23316 omhändertagandet 1
23317 omintetgör 2
23318 omintetgöra 1
23319 omintetgörs 1
23320 omistlig 1
23321 omkommit 1
23322 omkostnader 1
23323 omkostnadstäckning 4
23324 omkostnadstäckningen 1
23325 omkramad 1
23326 omkring 86
23327 omkringliggande 1
23328 omkull 1
23329 omkullkastar 1
23330 omlastning 1
23331 omlokaliseringar 3
23332 omlopp 9
23333 omloppsbana 1
23334 ommöblering 1
23335 omnämnande 1
23336 omnämnandena 1
23337 omnämnandet 1
23338 omnämnda 1
23339 omnämnde 1
23340 omnämns 2
23341 omoderna 1
23342 omodernt 2
23343 omogna 1
23344 omoralisk 1
23345 omoraliska 1
23346 omoraliskt 1
23347 omorganisation 1
23348 omorganisationen 7
23349 omorganisera 3
23350 omorganiserar 1
23351 omorganiseras 1
23352 omorganisering 1
23353 omorganiseringen 1
23354 omorientera 1
23355 omotiverat 2
23356 omplacera 1
23357 omplantering 1
23358 omprioritering 1
23359 ompröva 4
23360 omprövar 1
23361 omprövas 2
23362 omprövning 4
23363 omringades 1
23364 område 262
23365 områden 270
23366 områdena 56
23367 områdes 1
23368 områdesbegränsning 1
23369 områdesplaneringen 1
23370 området 221
23371 områdets 1
23372 omröstning 38
23373 omröstningar 9
23374 omröstningarna 5
23375 omröstningen 65
23376 omröstningen.1 1
23377 omröstningsförfarandet 1
23378 omröstningslistan 1
23379 omröstningsregistreringen 1
23380 omröstningsresultaten 1
23381 omsatts 1
23382 omsider 2
23383 omskolning 3
23384 omskrivningar 1
23385 omskärelsen 1
23386 omslag 1
23387 omslaget 1
23388 omsorg 16
23389 omsorgsfulla 1
23390 omsorgsfullt 5
23391 omstridd 3
23392 omstridda 1
23393 omstritt 2
23394 omstrukturera 4
23395 omstrukturering 20
23396 omstruktureringar 7
23397 omstruktureringarna 3
23398 omstruktureringen 2
23399 omstrukturerings- 1
23400 omstruktureringsplan 2
23401 omstruktureringsplaner 1
23402 omstuvning 1
23403 omställningar 1
23404 omställningen 1
23405 omställningsfasen 1
23406 omständighet 5
23407 omständigheten 3
23408 omständigheter 62
23409 omständigheterna 8
23410 omständliga 2
23411 omsvep 3
23412 omsvängning 2
23413 omsätta 8
23414 omsättas 4
23415 omsätter 1
23416 omsättning 3
23417 omsätts 4
23418 omtalade 4
23419 omtanke 1
23420 omtumlande 1
23421 omtvistad 1
23422 omtvistade 1
23423 omtvistat 1
23424 omvandla 3
23425 omvandlades 1
23426 omvandlas 4
23427 omvandlats 2
23428 omvandling 4
23429 omvandlingen 1
23430 omvandlingsprocess 1
23431 omvandlingsprocesser 1
23432 omväg 2
23433 omvägen 1
23434 omvälvande 1
23435 omvälvning 1
23436 omvälvningar 2
23437 omvänd 3
23438 omvända 4
23439 omvänt 7
23440 omvärdera 4
23441 omvärderas 2
23442 omvärdering 2
23443 omvärderingsperioden 1
23444 omvärld 1
23445 omvärlden 2
23446 omväxlande 2
23447 omvårdnad 1
23448 omänsklig 2
23449 omärkliga 1
23450 omärkligt 1
23451 omätliga 1
23452 omöjlig 5
23453 omöjliga 6
23454 omöjligen 2
23455 omöjliggjorde 1
23456 omöjliggör 1
23457 omöjliggörs 2
23458 omöjlighet 1
23459 omöjligheten 1
23460 omöjligt 27
23461 on 2
23462 ond 1
23463 onda 6
23464 ondo 2
23465 ondska 1
23466 ondskan 1
23467 ondskefulla 2
23468 ondskefullt 1
23469 one-stop-shop 1
23470 onekligen 4
23471 online-avtal 1
23472 online-ekonomin 1
23473 onsdag 7
23474 onsdagen 5
23475 onsdags 1
23476 ont 7
23477 onyanserat 1
23478 onödan 1
23479 onödig 6
23480 onödiga 7
23481 onödigt 9
23482 oomkullrunkeliga 1
23483 oomtvistad 1
23484 oordnad 1
23485 oordningen 2
23486 opaler 1
23487 opartisk 1
23488 opartiskhet 1
23489 opartiskt 4
23490 operahus 1
23491 operan 1
23492 operation 2
23493 operationer 4
23494 operativ 2
23495 operativa 9
23496 operativt 4
23497 operators 1
23498 operatör 1
23499 operatörer 1
23500 operatörerna 2
23501 operera 1
23502 opersonliga 1
23503 opinion 6
23504 opinionen 13
23505 opinioner 2
23506 opinionsbildare 1
23507 opinionsundersökningar 1
23508 oportunidades 1
23509 opp 5
23510 oppe 2
23511 opponera 3
23512 opportunism 1
23513 opportunister 1
23514 opposition 5
23515 oppositionell 1
23516 oppositionen 4
23517 oppositionens 2
23518 oppositionsledaren 1
23519 oppositionspolitikern 1
23520 oppositionstidningar 1
23521 opraktiskt 2
23522 oproportionerliga 2
23523 oproportionerligt 2
23524 optimal 4
23525 optimala 2
23526 optimalt 4
23527 optimera 1
23528 optimeras 1
23529 optimeringen 1
23530 optimism 5
23531 optimistisk 5
23532 optimistiska 2
23533 optimistiskt 4
23534 optioner 3
23535 optionskontrakt 1
23536 optiskt 1
23537 opålitlig 1
23538 orakel 1
23539 orange 1
23540 ord 166
23541 orda 4
23542 ordalag 13
23543 ordalydelsen 2
23544 ordats 1
23545 orden 21
23546 ordentlig 13
23547 ordentliga 1
23548 ordentligt 25
23549 order 4
23550 orders 1
23551 ordet 58
23552 ordförande 202
23553 ordförandebänken 1
23554 ordförandekolleger 1
23555 ordförandeland 1
23556 ordförandelandet 3
23557 ordföranden 25
23558 ordförandena 6
23559 ordförandens 3
23560 ordförandes 1
23561 ordförandeskap 44
23562 ordförandeskapen 2
23563 ordförandeskapens 1
23564 ordförandeskapet 120
23565 ordförandeskapets 31
23566 ordförandeskaps 3
23567 ordförandeskapsprogram 1
23568 ordförandestaten 1
23569 ordinarie 1
23570 ordinär 1
23571 ordlista 1
23572 ordna 6
23573 ordnade 3
23574 ordnandet 1
23575 ordnar 2
23576 ordnas 1
23577 ordnat 2
23578 ordnats 1
23579 ordning 28
23580 ordningar 1
23581 ordningen 13
23582 ordningsfråga 11
23583 ordningsfrågor 2
23584 ordningsfrågorna 2
23585 ordningsföljden 1
23586 ordningsmakt 1
23587 ordre 1
23588 ordrikt 2
23589 ordspråk 1
23590 ordspråket 2
23591 ordvalet 2
23592 ordvrängare 1
23593 ordvändning 1
23594 ordväxlingen 1
23595 orealistisk 2
23596 orealistiska 4
23597 orealistiskt 6
23598 oreda 2
23599 oredan 1
23600 oredlighet 1
23601 oreflekterat 1
23602 oregelbundet 1
23603 oreglerade 1
23604 oreglerat 1
23605 organ 49
23606 organen 12
23607 organens 2
23608 organet 3
23609 organisation 25
23610 organisationen 14
23611 organisationens 1
23612 organisationer 63
23613 organisationerna 20
23614 organisationernas 4
23615 organisationers 2
23616 organisations 1
23617 organisationsgraden 1
23618 organisationskapacitet 1
23619 organisationsschema 1
23620 organisationsstruktur 1
23621 organisatoriska 3
23622 organisatoriskt 1
23623 organisera 19
23624 organiserad 4
23625 organiserade 11
23626 organiserades 2
23627 organiserar 6
23628 organiseras 7
23629 organiserats 1
23630 organisering 1
23631 organiskt 1
23632 organism 1
23633 organismer 24
23634 organs 1
23635 orientaliska 1
23636 orienten 1
23637 orienterad 2
23638 orienterar 1
23639 orienteras 1
23640 orientering 2
23641 orienteringen 1
23642 orienteringsprogrammen 1
23643 originalitet 2
23644 originalspråket 1
23645 originalversionen 3
23646 originella 4
23647 originellt 2
23648 oriktiga 6
23649 oriktigheter 1
23650 oriktigt 2
23651 orimlig 2
23652 orimliga 6
23653 orimligt 3
23654 orkade 2
23655 orkan 1
23656 orkanen 1
23657 orkaner 1
23658 orkester 1
23659 orkestrarnas 1
23660 orm 4
23661 ormen 1
23662 ormens 2
23663 oro 100
23664 oroa 6
23665 oroad 6
23666 oroade 10
23667 oroande 23
23668 oroar 20
23669 oroas 1
23670 orolig 9
23671 oroliga 13
23672 oroligheter 1
23673 oron 17
23674 orosmoln 2
23675 orosmoment 5
23676 oroväckande 6
23677 orsak 11
23678 orsak-verkanrelationen 1
23679 orsaka 9
23680 orsakade 7
23681 orsakar 10
23682 orsakas 6
23683 orsakat 9
23684 orsakats 7
23685 orsaken 14
23686 orsaker 13
23687 orsakerna 12
23688 orsakssamband 1
23689 ort 4
23690 orten 3
23691 orter 2
23692 orthomixomicrovirus 1
23693 ortodoxa 1
23694 orubblig 2
23695 orubbliga 2
23696 orwellskt 1
23697 oräkneliga 2
23698 oräkneligt 1
23699 orätt 4
23700 orättfärdiga 1
23701 orättfärdigt 1
23702 orättvis 5
23703 orättvisa 4
23704 orättvisor 7
23705 orättvisorna 3
23706 orättvist 5
23707 orörda 1
23708 orörlig 3
23709 orörlighet 1
23710 orörligt 1
23711 osagt 1
23712 osammanhängande 4
23713 osanna 2
23714 osannolika 3
23715 osar 1
23716 osjälvisk 1
23717 osjälvständiga 1
23718 oskadliga 2
23719 oskarpa 1
23720 oskiljaktig 1
23721 oskiljaktiga 1
23722 oskriven 1
23723 oskuld 1
23724 oskuldsfull 1
23725 oskuldsfullt 1
23726 oskyldig 2
23727 oskyldiga 2
23728 oskyldigt 1
23729 oslipad 1
23730 osmidig 1
23731 osmältbar 1
23732 osolidariskt 1
23733 oss 1017
23734 ost 2
23735 ostraffade 1
23736 ostron 1
23737 ostronanläggningarna 1
23738 ostronodlare 3
23739 ostronodlarna 2
23740 ostronodling 1
23741 ostronodlingarna 1
23742 ostronodlingarnas 1
23743 ostronodlingen 1
23744 ostrukturerade 1
23745 ostört 1
23746 osv 3
23747 osv. 25
23748 osynlig 2
23749 osynliga 1
23750 osynligt 2
23751 osystematiskt 1
23752 osäker 2
23753 osäkerhet 18
23754 osäkerheten 2
23755 osäkert 2
23756 osäkra 5
23757 osäkrad 1
23758 osäkrare 1
23759 osårbart 1
23760 otacksamma 1
23761 otaliga 3
23762 otillfredsställande 3
23763 otillgängliga 1
23764 otillräcklig 10
23765 otillräckliga 12
23766 otillräcklighet 3
23767 otillräckligheten 1
23768 otillräckligt 10
23769 otillständigt 1
23770 otillåtliga 1
23771 otillåtligt 3
23772 otillåtna 1
23773 otjänst 2
23774 otrevligt 1
23775 otrolig 1
23776 otroliga 2
23777 otroligt 3
23778 otrygga 2
23779 otrygghet 1
23780 otryggt 1
23781 otvetydiga 4
23782 otvetydigt 2
23783 otvivelaktig 1
23784 otvivelaktigt 11
23785 otydlig 6
23786 otydliga 3
23787 otydlighet 1
23788 otydligt 4
23789 otyglad 2
23790 otympligt 1
23791 otäckheter 1
23792 otäckt 1
23793 otänkbart 5
23794 otålig 2
23795 otåliga 1
23796 otålighet 2
23797 otåligt 1
23798 ou 2
23799 oumbärlig 2
23800 oumbärliga 2
23801 oumbärligt 4
23802 oundgänglig 1
23803 oundgängliga 4
23804 oundgängligt 1
23805 oundviklig 1
23806 oundvikliga 9
23807 oundvikligen 5
23808 oundvikligt 5
23809 oupphörlig 1
23810 oupphörliga 2
23811 oupplösligt 1
23812 ouppmärksam 1
23813 outbildade 1
23814 outgrundlig 1
23815 outgrundligt 1
23816 outhärdlig 1
23817 outhärdliga 2
23818 outhärdligt 1
23819 outnyttjad 1
23820 outnyttjade 2
23821 outsinlig 1
23822 outsourcing 1
23823 outtalad 1
23824 outtömlig 1
23825 outtömligt 1
23826 ovala 1
23827 ovan 5
23828 ovana 1
23829 ovanför 7
23830 ovanifrån 2
23831 ovanlig 2
23832 ovanliga 3
23833 ovanligt 8
23834 ovannämnda 5
23835 ovanpå 5
23836 ovanstående 3
23837 ovederhäftigt 1
23838 over 2
23839 overall 2
23840 overhead-kostnader 1
23841 overkliga 1
23842 overkligt 1
23843 overksam 1
23844 overksamma 1
23845 ovetande 2
23846 oviktigt 1
23847 ovilja 3
23848 ovillkorligen 2
23849 ovisshet 1
23850 oväder 2
23851 ovädren 1
23852 ovädret 1
23853 oväld 1
23854 ovälkomna 1
23855 oväntade 3
23856 oväntat 5
23857 ovärderlig 2
23858 ovärdig 1
23859 ovärdiga 3
23860 ovärdigt 1
23861 oväsen 1
23862 oväsentligt 1
23863 oändlig 3
23864 oändliga 2
23865 oändlighet 3
23866 oändligt 3
23867 oåterkallelig 1
23868 oönskad 2
23869 oönskade 4
23870 oöverlagt 1
23871 oöverskådligt 1
23872 oöverstiglig 3
23873 oöverstigligt 1
23874 oövervinneligt 1
23875 p.17 1
23876 p.g.a. 4
23877 packa 3
23878 packad 1
23879 packat 2
23880 padanska 1
23881 paddlades 1
23882 paket 6
23883 paketet 3
23884 paketsektorn 1
23885 pakten 1
23886 palatsgrindarna 1
23887 palestinier 3
23888 palestinierna 8
23889 palestinsk 2
23890 palestinska 22
23891 palestinskt 2
23892 pallen 1
23893 pampig 1
23894 pandemiska 1
23895 paneler 2
23896 panelerna 1
23897 panga 1
23898 panik 3
23899 panikspridning 1
23900 panna 1
23901 pannan 4
23902 pannor 1
23903 panorama 2
23904 pansarvagnar 1
23905 pantomimiskt 1
23906 papegoja 1
23907 papp 3
23908 pappa 5
23909 papper 9
23910 papperet 3
23911 pappersarbete 4
23912 pappersarbetet 2
23913 pappersdokument 1
23914 papperskorgen 1
23915 pappersluntor 1
23916 pappersplaner 1
23917 papperstigrar 1
23918 pappersvaror 1
23919 par 50
23920 paradigm 3
23921 paradigmskifte 1
23922 paradis 1
23923 paradox 3
23924 paradoxal 3
23925 paradoxala 2
23926 paradoxalt 2
23927 paragrafrytteriet 1
23928 parallella 9
23929 parallellt 9
23930 paralyseras 1
23931 parameter 1
23932 parametern 1
23933 parametrar 1
23934 parametrarna 1
23935 paramilitära 1
23936 paramilitärt 1
23937 paraply 1
23938 paras 1
23939 parasiter 1
23940 parcours 1
23941 parece 2
23942 parentes 1
23943 paret 2
23944 parfym 1
23945 paria 1
23946 paritet 1
23947 parité 1
23948 park 1
23949 parken 2
23950 parkens 1
23951 parker 2
23952 parkerad 1
23953 parkerade 2
23954 parkerar 1
23955 parkeringskort 2
23956 parkeringsplatser 1
23957 parlament 135
23958 parlamentariker 14
23959 parlamentarikerna 3
23960 parlamentarisk 11
23961 parlamentariska 18
23962 parlamentariskt 4
23963 parlamentarismen 1
23964 parlamenten 24
23965 parlamentens 2
23966 parlamentet 525
23967 parlamentet- 1
23968 parlamentets 127
23969 parlaments 5
23970 parlamentsbesluten 1
23971 parlamentsbyggnaden 1
23972 parlamentsdebatt 3
23973 parlamentsforum 1
23974 parlamentsgrupp 1
23975 parlamentskolleger 2
23976 parlamentskollegerna 1
23977 parlamentsledamot 16
23978 parlamentsledamoten 3
23979 parlamentsledamöter 29
23980 parlamentsledamöterna 9
23981 parlamentsledamöternas 1
23982 parlamentsnivå 1
23983 parlamentspresidiets 1
23984 parlamentsutskott 3
23985 parlamentsutskotten 1
23986 parlamentsutskottet 1
23987 parmaskinkstunga 1
23988 parningsplatser 1
23989 parodi 1
23990 part 9
23991 parten 3
23992 parter 50
23993 parterna 16
23994 parternas 11
23995 parters 4
23996 parti 49
23997 partiapparaterna 1
23998 partiell 1
23999 partiella 3
24000 partier 24
24001 partierna 13
24002 partiernas 5
24003 partiers 2
24004 partiet 18
24005 partiets 29
24006 partigrupp 3
24007 partigruppen 1
24008 partiintressen 1
24009 partikrati 1
24010 partiledare 1
24011 partimedlems 1
24012 partipolitisk 1
24013 partipolitiska 2
24014 partiprogram 3
24015 partiprogrammet 1
24016 partis 3
24017 partisk 1
24018 partiska 2
24019 partiskt 1
24020 partisplittringens 1
24021 partivänner 1
24022 partner 31
24023 partnern 1
24024 partnerparti 1
24025 partnerrelationen 1
24026 partners 4
24027 partnership 1
24028 partnerskap 41
24029 partnerskapen 3
24030 partnerskapens 1
24031 partnerskapet 8
24032 partnerskapets 2
24033 partnerskaps- 1
24034 partnerskapsavtal 4
24035 partnerskapsavtalen 1
24036 partnerskapsavtalet 4
24037 partnerskapsbidrag 1
24038 partnerskapsformer 1
24039 partnerskapskonceptet 1
24040 partnerskapsländerna 1
24041 partnerskapsmålet 1
24042 partnerskapspolitiken 1
24043 partnerskapsprincipen 3
24044 partnerskapsrådet 1
24045 partnerskapsuppgörelserna 1
24046 partnerstater 1
24047 parts 1
24048 party 1
24049 partyt 1
24050 pas 2
24051 pass 10
24052 passa 10
24053 passade 3
24054 passadvind 1
24055 passage 2
24056 passagerarbuss 1
24057 passagerare 5
24058 passagerarna 6
24059 passagerarnas 1
24060 passagerartransporter 1
24061 passande 10
24062 passar 12
24063 passera 5
24064 passerade 4
24065 passerar 1
24066 passerat 2
24067 passet 1
24068 passion 3
24069 passionerat 1
24070 passiv 1
24071 passivitet 1
24072 passiviteten 1
24073 passivt 2
24074 passusen 1
24075 pastellmjuka 1
24076 patent 5
24077 patentfrågorna 1
24078 patentmediciner 1
24079 patenträtt 1
24080 patenträttigheterna 1
24081 patentslag 1
24082 paternalistiska 2
24083 paternalistiskt 1
24084 patetisk 1
24085 patetiskt 1
24086 patient 1
24087 patienter 3
24088 patogen 1
24089 patologiska 1
24090 patriarkalisk 1
24091 patriot 1
24092 patrioters 1
24093 patriotism 1
24094 patrullbåt 1
24095 paus 4
24096 pausen 1
24097 pauser 1
24098 paying 1
24099 peanuts-belopp 1
24100 pedagogiska 2
24101 pedagogiskt 1
24102 pedofilskandaler 1
24103 peka 17
24104 pekade 10
24105 pekar 16
24106 pekat 9
24107 pelare 10
24108 pelaren 8
24109 pelarna 7
24110 pengar 94
24111 pengarna 31
24112 penndrag 1
24113 penning- 1
24114 penningdyrkan 1
24115 penningflöden 1
24116 penningflödena 1
24117 penningfurstars 1
24118 penninggirig 1
24119 penningmarknad 1
24120 penningmarknadsinstrument 1
24121 penningmedel 1
24122 penningpolitik 3
24123 penningpolitiken 2
24124 penningpolitisk 1
24125 penningpolitiska 3
24126 penningreferenser 1
24127 penningresurser 1
24128 penningstabilitet 1
24129 penningsummor 1
24130 penningtvätt 4
24131 penningväsendets 1
24132 pension 8
24133 pensioner 10
24134 pensioneras 1
24135 pensionerna 8
24136 pensionsbomben 1
24137 pensionsfonder 5
24138 pensionsfondernas 1
24139 pensionsförmånerna 1
24140 pensionsförsäkringarna 1
24141 pensionsmedlen 1
24142 pensionspolitik 1
24143 pensionsrättigheter 1
24144 pensionssystem 2
24145 pensionssystemen 3
24146 pensionssystemens 1
24147 pensionssystemet 2
24148 pensionstidbomb 1
24149 pensionär 3
24150 pensionärer 3
24151 pensionärerna 1
24152 pensionärernas 1
24153 pensionärers 1
24154 per 60
24155 perfekt 11
24156 perfekta 2
24157 pergamentrulle 1
24158 perifera 10
24159 periferin 2
24160 perifert 1
24161 period 32
24162 perioden 60
24163 perioder 5
24164 perioderna 2
24165 periodisk 1
24166 periodiska 15
24167 periodvis 1
24168 perito 1
24169 permanent 7
24170 permanenta 6
24171 perrongen 1
24172 person 32
24173 persona 2
24174 personal 29
24175 personalbrist 1
24176 personaldelen 1
24177 personalen 4
24178 personalens 1
24179 personalförstärkning 1
24180 personalnedskärningar 2
24181 personalnedskärningarna 1
24182 personalpolitik 3
24183 personalpolitiken 1
24184 personalresurser 2
24185 personalresurserna 2
24186 personalsidan 1
24187 personalstrukturen 1
24188 personalutbildning 2
24189 personbil 1
24190 personbyte 1
24191 personell 1
24192 personella 2
24193 personen 2
24194 personer 128
24195 personerna 7
24196 personernas 1
24197 personers 6
24198 personifieras 1
24199 personlandminor 3
24200 personlig 5
24201 personliga 24
24202 personligen 33
24203 personlighet 1
24204 personligheten 1
24205 personligt 4
24206 personne 1
24207 persons 2
24208 persontransporter 1
24209 perspektiv 45
24210 perspektivet 7
24211 peruaner 1
24212 perversas 1
24213 pessimistisk 1
24214 pessimistiskt 1
24215 pesten 3
24216 pestens 1
24217 petar 1
24218 petition 1
24219 petroleum 1
24220 pharmaceutiques 1
24221 phtalater 1
24222 pickade 1
24223 pickar 1
24224 pickelsburk 1
24225 pickles 1
24226 picknickväska 1
24227 pigg 1
24228 pikade 1
24229 pil 1
24230 pilgrimer 2
24231 pilgrimerna 1
24232 piloten 1
24233 piloter 1
24234 pilotfunktion 1
24235 pilotmervärde 1
24236 pilotprogram 2
24237 pilotprojekt 14
24238 pilotstudier 1
24239 pincene 1
24240 pinglade 1
24241 pinsam 2
24242 pinsamt 2
24243 pionjärer 1
24244 pionjärerna 1
24245 pip 1
24246 pipa 1
24247 pipande 1
24248 pipor 1
24249 pipskägg 1
24250 pir 1
24251 pirat 1
24252 pirater 2
24253 piraternas 1
24254 piratkopiering 1
24255 piratkopior 1
24256 piratversion 1
24257 pirerna 1
24258 pivotabellvy 2
24259 pivotdiagramkomponenten 1
24260 pivotdiagramvy 2
24261 pivotdiagramvyns 1
24262 pivottabell 2
24263 pivottabell- 1
24264 pivottabellen 2
24265 pivottabellens 1
24266 pivottabeller 2
24267 pivottabellista 7
24268 pivottabellistan 1
24269 pivottabellistans 1
24270 pivottabellistor 2
24271 pivottabellkomponenten 2
24272 pivottabellvy 5
24273 pivottabellvyer 3
24274 pivottabellvyn 5
24275 pivottabellvyns 1
24276 pivottabelläge 2
24277 pivottabelläget 2
24278 pjäser 1
24279 placera 12
24280 placerad 4
24281 placerade 3
24282 placerades 2
24283 placerar 8
24284 placeras 8
24285 placerat 5
24286 placerats 1
24287 placering 2
24288 placeringen 1
24289 placeringsformerna 1
24290 placeringsmarknaden 2
24291 placeringsmöjligheterna 1
24292 pladask 1
24293 pladder 1
24294 plagg 1
24295 plan 41
24296 planekonomiska 1
24297 planen 9
24298 planens 1
24299 planer 32
24300 planera 8
24301 planerad 5
24302 planerade 24
24303 planerades 3
24304 planerande 1
24305 planerar 24
24306 planeras 13
24307 planerat 8
24308 planerats 4
24309 planering 24
24310 planeringen 12
24311 planeringsfasen 2
24312 planeringsskedet 2
24313 planeringsstadiet 1
24314 planerna 7
24315 planet 34
24316 planeten 3
24317 planetens 2
24318 planeter 3
24319 planets 2
24320 plankton 1
24321 planlagda 1
24322 planläggning 1
24323 planlösa 2
24324 planlösningen 1
24325 planlöst 2
24326 plantera 1
24327 plantor 1
24328 plast 6
24329 plastbagar 1
24330 plastdisk 1
24331 plasten 1
24332 plastväv 1
24333 plats 82
24334 platsen 17
24335 platser 32
24336 platserna 3
24337 platt 2
24338 platta 3
24339 plattades 1
24340 plattan 2
24341 plattare 1
24342 plattform 1
24343 plattformar 1
24344 plattheter 1
24345 playing 1
24346 plenardebatten 1
24347 plenarkammaren 2
24348 plenarsalen 1
24349 plenarsammanträde 4
24350 plenarsammanträden 1
24351 plenarsammanträdena 1
24352 plenarsammanträdet 7
24353 plenisalen 2
24354 plenum 9
24355 plenumet 2
24356 plikt 11
24357 plikten 2
24358 pliktskyldig 1
24359 plimsollmärket 1
24360 plocka 4
24361 plockade 3
24362 plockats 1
24363 plumpa 1
24364 plundra 2
24365 plundrare 1
24366 plundras 1
24367 plundring 1
24368 plundringarna 1
24369 plundringen 1
24370 pluralism 1
24371 pluralistiska 4
24372 pluralistiskt 1
24373 plus 5
24374 pluskonto 1
24375 plädera 2
24376 pläderar 5
24377 pläderingen 1
24378 plätt 1
24379 plåga 1
24380 plågade 2
24381 plågar 1
24382 plågas 1
24383 plånboken 1
24384 plånböcker 1
24385 plåt 2
24386 plåtdunk 1
24387 plåtskjul 1
24388 plötslig 3
24389 plötsliga 1
24390 plötsligt 37
24391 poche 1
24392 poena 1
24393 poet 4
24394 poetromantiska 1
24395 pojkar 2
24396 pojkarna 1
24397 pojke 10
24398 pojken 8
24399 pojkes 1
24400 polacker 1
24401 polariserat 1
24402 poldermodellen 1
24403 pole 1
24404 polemik 2
24405 polemisk 1
24406 polemiskt 1
24407 polera 1
24408 policy 7
24409 policybeslut 1
24410 policydel 1
24411 policyförslag 1
24412 policyn 2
24413 policyutveckling 1
24414 polis 7
24415 polis- 1
24416 polisakademi 1
24417 polisbevakning 3
24418 polisbyrån 1
24419 polisen 13
24420 polisenheter 1
24421 polisens 1
24422 poliser 16
24423 polisexperter 1
24424 polisfrågan 1
24425 polisiär 2
24426 polisiära 7
24427 poliskommissarien 1
24428 poliskåren 1
24429 polismyndigheterna 2
24430 polissamarbetet 1
24431 polisstyre 1
24432 polisstyrka 2
24433 polisstyrkan 2
24434 polisstyrkor 1
24435 polisstyrkorna 1
24436 polistjänstemän 2
24437 polisväsendet 1
24438 political 1
24439 politik 314
24440 politiken 110
24441 politikens 7
24442 politiker 27
24443 politikerjargong 1
24444 politikerna 1
24445 politikernas 1
24446 politikers 1
24447 politikområde 4
24448 politikområden 51
24449 politikområdena 6
24450 politikområdenas 2
24451 politiks 2
24452 politiseras 1
24453 politiserat 1
24454 politisk 121
24455 politisk-ekonomiska 1
24456 politiska 374
24457 politiskt 87
24458 polsk 2
24459 polska 3
24460 polske 1
24461 polyaromatisk 1
24462 polycentrisk 1
24463 pompöst 1
24464 pool 1
24465 popularisera 1
24466 populism 1
24467 populismen 1
24468 populistisk 1
24469 populistiska 2
24470 populära 3
24471 porslin 1
24472 porslinsbutik 1
24473 port 1
24474 port-state 2
24475 porten 3
24476 portfölj 4
24477 portföljen 1
24478 portföljer 2
24479 portföljförvaltning 1
24480 portmonnäer 1
24481 portmonnän 1
24482 portokostnad 1
24483 porttelefonen 1
24484 portugis 1
24485 portugisisk 3
24486 portugisiska 126
24487 portugisiske 5
24488 portugisiskt 3
24489 portvin 2
24490 posidonia 1
24491 position 10
24492 positionen 3
24493 positioner 6
24494 positiv 68
24495 positiva 72
24496 positivlista 3
24497 positivlistan 1
24498 positivt 81
24499 post 9
24500 posta 1
24501 postala 1
24502 postanställdas 2
24503 postavgifterna 1
24504 postbefordran 1
24505 postbrevbärarna 1
24506 postdirektivet 2
24507 postdistribuerad 1
24508 posten 23
24509 postens 2
24510 poster 11
24511 posterna 4
24512 postföretag 1
24513 postföretagen 4
24514 postförsändelsernas 1
24515 postgången 1
24516 posthandeln 1
24517 posthanteringen 1
24518 postindustriell 1
24519 postindustriella 1
24520 postkoloniala 1
24521 postkontor 13
24522 postkontoren 7
24523 postkontorens 1
24524 postkontoret 2
24525 postkontorsnätverket 1
24526 postkontorstjänster 1
24527 postlåda 1
24528 postmannen 1
24529 postmarknaden 4
24530 postmilitär 1
24531 postmonopolet 1
24532 postområdet 1
24533 postoperatörer 1
24534 postoperatörerna 2
24535 postpolitiken 1
24536 postsektorn 6
24537 postsektorns 2
24538 postservice 2
24539 postsystem 1
24540 posttjänst 2
24541 posttjänstdirektivet 3
24542 posttjänsten 3
24543 posttjänstens 1
24544 posttjänster 29
24545 posttjänsterna 30
24546 posttjänstesektorn 1
24547 posttrafiken 1
24548 postturer 1
24549 posttömningen 1
24550 postutbärare 1
24551 postutbärning 1
24552 postutdelning 2
24553 postutställd 1
24554 postverk 2
24555 postverken 4
24556 postverket 3
24557 postverkets 1
24558 postverksamheten 1
24559 postväsendet 4
24560 potatis 1
24561 potential 13
24562 potentialen 1
24563 potentialer 1
24564 potentiell 3
24565 potentiella 12
24566 potentiellt 3
24567 pottaska 1
24568 poäng 3
24569 poängen 1
24570 poängsystem 4
24571 poängtera 11
24572 poängterar 4
24573 poängterat 3
24574 poängterats 1
24575 ppm 1
24576 prackats 1
24577 practice 1
24578 practice-metoder 1
24579 practices 2
24580 pragmatisk 2
24581 pragmatiska 2
24582 pragmatiskt 2
24583 pragmatism 1
24584 praktexempel 1
24585 praktfull 1
24586 praktfullt 1
24587 praktik 3
24588 praktikanter 2
24589 praktiken 35
24590 praktiserar 1
24591 praktiseras 1
24592 praktisk 9
24593 praktiska 33
24594 praktiskt 23
24595 prat 3
24596 prata 14
24597 pratade 1
24598 pratar 3
24599 pratat 2
24600 pratet 1
24601 praxis 14
24602 praxisen 1
24603 precedensfall 1
24604 precis 93
24605 precisa 5
24606 precisera 5
24607 preciserad 1
24608 preciserade 2
24609 preciserar 3
24610 preciseras 2
24611 preciserat 1
24612 precisering 3
24613 preciseringar 5
24614 precision 5
24615 precist 1
24616 predika 1
24617 predikande 1
24618 prefekt 1
24619 prefektemblem 1
24620 prefekts 1
24621 preferens 2
24622 preferensbehandla 1
24623 preferenser 3
24624 preferensoptionen 1
24625 preferenssystemet 2
24626 prejudicerande 1
24627 prejudikat 5
24628 preliminära 5
24629 preliminärt 1
24630 premiss 1
24631 premisser 1
24632 premisserna 1
24633 premiärminister 22
24634 premiärministern 9
24635 premiärministrar 1
24636 premiärministrarna 1
24637 prerogativ 4
24638 prerogativet 1
24639 present 4
24640 presentabla 1
24641 presentation 5
24642 presentationen 4
24643 presentations- 1
24644 presentationsfilen 1
24645 presentationsformat 3
24646 presentationsinformation 1
24647 presentationsinformationen 1
24648 presenter 3
24649 presentera 21
24650 presenterade 7
24651 presenterades 5
24652 presenterandet 1
24653 presenterar 7
24654 presenteras 12
24655 presenterat 7
24656 presenterats 2
24657 president 29
24658 presidenten 8
24659 presidentens 1
24660 presidenter 1
24661 presidentestraden 1
24662 presidentvalet 1
24663 presidiet 4
24664 presidiets 1
24665 presidium 1
24666 press 8
24667 pressa 3
24668 pressade 5
24669 pressande 1
24670 pressar 2
24671 pressen 15
24672 pressens 2
24673 pressfotografer 1
24674 pressfrihet 5
24675 pressfriheten 2
24676 presskonferens 1
24677 presskonferenser 2
24678 pressmeddelande 1
24679 pressorgan 1
24680 presstjänst 1
24681 prestanda 3
24682 prestation 5
24683 prestationer 2
24684 prestationerna 1
24685 prestationsförmågan 2
24686 prestera 2
24687 presterat 1
24688 preventiv 1
24689 preventiva 1
24690 preventivt 1
24691 prick 1
24692 pricka 1
24693 prickar 1
24694 prickfritt 1
24695 prima 1
24696 primitiva 2
24697 primära 2
24698 primärsektorernas 1
24699 primärt 2
24700 princip 73
24701 principen 98
24702 principer 78
24703 principerna 33
24704 principernas 1
24705 principfast 1
24706 principfrågor 2
24707 principförklaring 1
24708 principförklaringar 1
24709 principiell 1
24710 principiella 3
24711 principiellt 14
24712 principskäl 1
24713 principöverenskommelse 1
24714 prinsessan 1
24715 priori 4
24716 prioritera 21
24717 prioriterad 5
24718 prioriterade 16
24719 prioriterades 1
24720 prioriterar 9
24721 prioriteras 16
24722 prioriterat 5
24723 prioritering 7
24724 prioriteringar 31
24725 prioriteringarna 9
24726 prioriteringen 7
24727 prioriteringslistan 1
24728 prioriteringsområden 1
24729 prioriteringsskala 1
24730 prioritet 12
24731 prioriteter 7
24732 prioriteterna 4
24733 priorssäte 1
24734 pris 25
24735 pris- 2
24736 prisa 1
24737 prisas 1
24738 prisats 1
24739 prisberäkningar 1
24740 priser 16
24741 priserna 12
24742 priset 24
24743 prisfastställandet 1
24744 prisgränser 1
24745 prisgränserna 2
24746 prishöjningar 1
24747 prisnivåerna 1
24748 prispolitik 1
24749 prispolitiken 3
24750 prisskillnader 1
24751 prisstabilitet 4
24752 prisstegring 1
24753 prissänkning 1
24754 prissänkningar 1
24755 prissättning 1
24756 prissättningen 2
24757 prisutvecklingen 1
24758 prisökning 2
24759 prisökningen 1
24760 privat 8
24761 privata 54
24762 privatekonomin 1
24763 privatiseras 1
24764 privatisering 9
24765 privatiseringar 2
24766 privatiseringarna 1
24767 privatiseringen 3
24768 privatiseringens 1
24769 privatlivet 1
24770 privatperson 1
24771 privatpersoner 2
24772 privatsfär 1
24773 privilege 2
24774 privilegier 3
24775 privilegiera 1
24776 privilegierade 2
24777 privilegiet 1
24778 privilegium 4
24779 priviligierade 1
24780 proaktiv 3
24781 problem 365
24782 problematik 1
24783 problematiken 5
24784 problematisk 2
24785 problematiska 1
24786 problematiskt 2
24787 problemen 70
24788 problemens 2
24789 problemet 117
24790 problemets 3
24791 problemlista 1
24792 problemområden 1
24793 problemområdena 3
24794 procedur 3
24795 proceduren 1
24796 procedurer 3
24797 procedurreglerna 1
24798 procent 276
24799 procentandel 2
24800 procentandelarna 1
24801 procenten 3
24802 procents 3
24803 procentsats 3
24804 procentsatsen 1
24805 procentsatser 2
24806 procentsiffror 1
24807 procenttal 3
24808 procenttalet 1
24809 procenttecken 1
24810 procentuellt 1
24811 process 62
24812 processen 47
24813 processens 1
24814 processer 15
24815 processerna 4
24816 processfrågor 2
24817 procession 1
24818 processregler 1
24819 processrättens 1
24820 processuell 1
24821 processuella 4
24822 procès 1
24823 producent 3
24824 producentansvar 3
24825 producentansvaret 3
24826 producenten 6
24827 producentens 2
24828 producenter 11
24829 producenterna 6
24830 producentländerna 1
24831 producera 8
24832 producerade 1
24833 producerar 4
24834 produceras 4
24835 producerat 3
24836 producerats 1
24837 produkt 18
24838 produkten 7
24839 produktens 1
24840 produkter 42
24841 produkterna 4
24842 produkternas 4
24843 produktinnovationer 1
24844 produktion 13
24845 produktionen 5
24846 produktioner 2
24847 produktionsanläggningar 1
24848 produktionsföretag 1
24849 produktionskedjan 1
24850 produktionskostnad 1
24851 produktionskostnaderna 2
24852 produktionsled 1
24853 produktionsmedlen 1
24854 produktionsmetod 1
24855 produktionsmetoder 1
24856 produktionsmodell 1
24857 produktionsnedgången 1
24858 produktionsprocessen 1
24859 produktionsresurser 1
24860 produktionssektor 1
24861 produktionssystem 1
24862 produktionsverksamhet 1
24863 produktiv 4
24864 produktiva 8
24865 produktivitet 6
24866 produktiviteten 6
24867 produktivitetsmarginaler 1
24868 produktivitetsstegring 1
24869 produktivitetsvinster 2
24870 produktivitetsvinsterna 1
24871 produktivt 3
24872 produkts 3
24873 professionalism 2
24874 professionell 1
24875 professionella 4
24876 professor 11
24877 profeten 1
24878 profil 3
24879 profilen 1
24880 profilera 1
24881 profilerad 1
24882 profilerat 1
24883 profiterar 1
24884 profylaktisk 1
24885 prognos 2
24886 prognoserna 1
24887 program 227
24888 programansvariga 1
24889 programdokument 1
24890 programförklaring 2
24891 programinitiativen 1
24892 programinriktning 1
24893 programmatiskt 2
24894 programmen 53
24895 programmeringsspråk 1
24896 programmet 89
24897 programmets 5
24898 programmässiga 2
24899 programmål 1
24900 programperioden 4
24901 programplanering 4
24902 programplaneringen 3
24903 programplaneringsdokument 1
24904 programplaneringsperiod 1
24905 programplaneringsperioden 7
24906 programpunkt 1
24907 programrundan 1
24908 programs 1
24909 programutformningen 1
24910 programvaror 2
24911 programverksamhet 1
24912 progressiv 4
24913 progressiva 1
24914 progressivt 2
24915 prohibition 2
24916 projekt 150
24917 projektadministration 2
24918 projekten 26
24919 projektens 4
24920 projektet 26
24921 projektets 1
24922 projektförslagen 1
24923 projektil 1
24924 projektledningen 2
24925 projektresultat 1
24926 projekts 3
24927 projektvalet 1
24928 proklamera 2
24929 promenad 2
24930 promenaden 1
24931 promenader 2
24932 promenera 2
24933 promenerade 2
24934 promille 1
24935 prompt 1
24936 pronazistiskt 1
24937 propaganda 9
24938 propagandakampanj 1
24939 propagandaskyltar 1
24940 propagera 1
24941 propagerat 2
24942 proportion 6
24943 proportionalitet 1
24944 proportionalitetsprincipen 1
24945 proportionalitetsprinciperna 1
24946 proportionella 1
24947 proportionellt 2
24948 proportioner 2
24949 proportionerliga 1
24950 proppar 1
24951 propuesta 2
24952 prosaiska 1
24953 prospekt 3
24954 prostituerade 2
24955 prostitution 2
24956 prostitutionen 1
24957 proteininnehåll 1
24958 proteinkornspåse 1
24959 protektionism 6
24960 protektionistisk 1
24961 protektionistiska 2
24962 protest 6
24963 protestaktioner 1
24964 protestanter 1
24965 protestantiska 2
24966 protestantiskt 1
24967 protesten 1
24968 protester 7
24969 protestera 2
24970 protesterade 3
24971 protesterar 5
24972 protesterat 2
24973 protestljuden 1
24974 protokoll 13
24975 protokollen 7
24976 protokollet 33
24977 prov 22
24978 prova 1
24979 provanställda 1
24980 provet 1
24981 provins 3
24982 provinsen 4
24983 provinser 1
24984 provinserna 1
24985 provisorisk 2
24986 provisoriska 4
24987 provkandidaterna 1
24988 provkarta 1
24989 provocerande 1
24990 provokation 1
24991 provokationer 1
24992 provunderlag 1
24993 prydd 1
24994 prydligt 1
24995 prydnadssak 1
24996 prygla 1
24997 pryglades 1
24998 prägel 4
24999 prägeln 2
25000 prägla 3
25001 präglad 5
25002 präglade 3
25003 präglades 1
25004 präglar 2
25005 präglas 7
25006 präglat 1
25007 präglats 3
25008 pråmarna 1
25009 préparez 1
25010 pröva 3
25011 prövade 2
25012 prövar 1
25013 prövas 3
25014 prövats 1
25015 prövning 6
25016 prövningar 3
25017 prövningarna 1
25018 prövoår 1
25019 pseudo- 1
25020 psykiska 1
25021 psykiskt 1
25022 psykologiska 2
25023 psykologiskt 1
25024 pubar 2
25025 public 1
25026 publicera 1
25027 publicerade 1
25028 publicerades 2
25029 publiceras 1
25030 publicering 1
25031 publicitet 1
25032 publik 2
25033 publiken 1
25034 puertoricansk 1
25035 puffade 1
25036 pulserar 1
25037 pulvret 1
25038 pumpas 4
25039 pund 7
25040 punga 1
25041 pungslagna 1
25042 punkt 224
25043 punkten 83
25044 punkter 99
25045 punkterna 16
25046 punktlig 1
25047 punktligt 1
25048 punkts 1
25049 punktskattepliktiga 1
25050 punktskatter 11
25051 punktskattesats 1
25052 punktskattesatser 1
25053 punktskattesatserna 1
25054 pures 1
25055 puritanska 1
25056 purpurröda 1
25057 pussel 2
25058 pusselbit 1
25059 pusslet 1
25060 putande 1
25061 putsade 2
25062 putsmedel 1
25063 putstrasa 1
25064 pyjamasbyxor 1
25065 pyjamasen 2
25066 pyramidisk 1
25067 pälsverk 1
25068 pärla 1
25069 pärlband 1
25070 pärlbroderier 1
25071 pärlor 1
25072 pärmen 1
25073 päron 1
25074 på 6240
25075 påbjuder 1
25076 påbjudet 1
25077 påbörja 4
25078 påbörjade 3
25079 påbörjades 3
25080 påbörjar 1
25081 påbörjas 3
25082 påbörjat 8
25083 påbörjats 3
25084 pådrag 1
25085 pådrivandet 1
25086 pådyvlas 1
25087 påfallande 3
25088 påfrestande 1
25089 påfrestning 2
25090 påfrestningar 1
25091 påfrestningarnas 1
25092 påfyllning 1
25093 påföljande 2
25094 påföljd 2
25095 påföljden 1
25096 påföljder 3
25097 påföljderna 2
25098 påförde 1
25099 pågick 7
25100 pågå 4
25101 pågående 23
25102 pågår 32
25103 pågått 3
25104 påkalla 1
25105 påkallar 1
25106 påkommen 1
25107 påkopplad 1
25108 pålagor 3
25109 pålitlig 3
25110 pålitliga 2
25111 pålitlighet 1
25112 pålitligt 1
25113 pålägga 1
25114 påläggas 1
25115 påminda 1
25116 påminde 7
25117 påminna 85
25118 påminnande 1
25119 påminnas 2
25120 påminnelse 2
25121 påminner 28
25122 påmint 3
25123 påpeka 58
25124 påpekade 22
25125 påpekades 2
25126 påpekande 8
25127 påpekanden 9
25128 påpekandet 1
25129 påpekar 17
25130 påpekas 5
25131 påpekat 29
25132 påpekats 8
25133 påsen 1
25134 påsk 1
25135 påskynda 7
25136 påskyndande 1
25137 påskyndar 1
25138 påskyndas 4
25139 påstod 1
25140 påstods 1
25141 påstridiga 1
25142 påstå 17
25143 påstådd 1
25144 påstående 6
25145 påståenden 3
25146 påståendena 1
25147 påståendet 3
25148 påstår 13
25149 påstås 6
25150 påståtts 2
25151 påstötning 1
25152 påta 1
25153 påtaglig 4
25154 påtagliga 7
25155 påtagligen 1
25156 påtagligt 6
25157 påtala 3
25158 påtalade 2
25159 påtalar 1
25160 påtalat 3
25161 påtalats 5
25162 påtryckning 1
25163 påtryckningar 19
25164 påtryckningarna 2
25165 påtryckningsgrupper 2
25166 påtryckningskampanj 1
25167 påtryckningsmedel 4
25168 påtryckningssanktioner 1
25169 påträffades 1
25170 påträffas 1
25171 påtvinga 3
25172 påtvingad 2
25173 påtvingade 2
25174 påtvingar 1
25175 påtvingas 2
25176 påtvingats 1
25177 påverka 27
25178 påverkade 1
25179 påverkan 13
25180 påverkar 39
25181 påverkas 17
25182 påverkat 5
25183 påverkats 8
25184 påvisades 1
25185 påvisar 2
25186 påvisas 1
25187 påvisat 4
25188 påvisats 1
25189 påvisbart 1
25190 qua 3
25191 quality 1
25192 que 1
25193 quidditch 1
25194 quidditchlag 1
25195 quo 3
25196 quota-hoping 1
25197 r 1
25198 rabatt 1
25199 rabatterna 1
25200 rabbi 1
25201 rabbin 1
25202 racerkvast 1
25203 rad 72
25204 rad- 4
25205 raden 4
25206 rader 5
25207 radera 1
25208 raderna 3
25209 radfält 2
25210 radikal 7
25211 radikala 10
25212 radikalernas 1
25213 radikalisering 1
25214 radikalt 9
25215 radio 1
25216 radio- 3
25217 radioaktiva 1
25218 radioaktivt 1
25219 radioamatörfrågan 1
25220 radioklassrum 1
25221 radiologiska 2
25222 radion 4
25223 radioutsändningar 1
25224 radområdet 1
25225 raffinaderier 2
25226 raffinaderiägarna 1
25227 raggiga 1
25228 raiden 2
25229 rak 4
25230 raka 8
25231 rakade 1
25232 rakblad 1
25233 raketanfall 1
25234 raketerna 1
25235 rakryggade 1
25236 raksträcka 1
25237 rakt 14
25238 ram 41
25239 ramar 9
25240 ramarna 6
25241 ramavtal 4
25242 ramavtalet 2
25243 rambeslut 17
25244 rambeslutet 5
25245 rambestämmelser 2
25246 ramdirektiv 10
25247 ramdirektivet 7
25248 ramen 173
25249 ramförslaget 3
25250 ramkonventionen 1
25251 ramlade 4
25252 ramlagstiftning 1
25253 ramlat 1
25254 rammar 1
25255 rampljus 1
25256 rampljuset 1
25257 ramprogram 4
25258 ramprogrammen 1
25259 ramprogrammet 10
25260 ramverk 2
25261 ramvillkor 3
25262 ramvillkoren 2
25263 randområde 1
25264 randområden 9
25265 randområdena 20
25266 randområdet 1
25267 randregioner 1
25268 rang 1
25269 rangordningen 1
25270 rann 3
25271 rannsakar 1
25272 rapid 2
25273 rapning 1
25274 rapphöna 1
25275 rappningen 1
25276 rapport 104
25277 rapport.xml 1
25278 rapporten 55
25279 rapportens 4
25280 rapporter 31
25281 rapportera 8
25282 rapporterade 1
25283 rapporterades 1
25284 rapporterar 1
25285 rapporteras 2
25286 rapporterat 2
25287 rapporterats 1
25288 rapportering 5
25289 rapporterna 6
25290 rapportsiffror 1
25291 ras 6
25292 rasade 2
25293 rasande 4
25294 rasat 1
25295 raser 1
25296 rasera 2
25297 raseri 1
25298 rashatet 1
25299 rasisistiska 1
25300 rasism 27
25301 rasismen 5
25302 rasist 1
25303 rasisterna 1
25304 rasistisk 3
25305 rasistiska 18
25306 rasistiskt 5
25307 raskt 2
25308 rasmässig 1
25309 rasslade 2
25310 rast 1
25311 rastillhörighet 1
25312 rastlös 1
25313 rastlösa 2
25314 ratar 1
25315 ratificera 2
25316 ratificerad 1
25317 ratificerade 1
25318 ratificerades 1
25319 ratificerar 4
25320 ratificeras 1
25321 ratificerat 7
25322 ratificerats 2
25323 ratificering 2
25324 ratificeringen 3
25325 ratificeringsförfarandet 1
25326 ratificeringshandlingar 1
25327 ratificeringsprocessen 2
25328 rating 2
25329 rationalisera 5
25330 rationaliserad 1
25331 rationaliserar 1
25332 rationalisering 3
25333 rationaliseringen 1
25334 rationaliseringseffekterna 1
25335 rationell 5
25336 rationella 2
25337 rationellt 5
25338 ratten 1
25339 ravin 1
25340 razzia 2
25341 razzior 1
25342 re-admission 1
25343 reaction 2
25344 reagera 24
25345 reagerade 2
25346 reagerar 7
25347 reagerat 4
25348 reaktion 16
25349 reaktioner 7
25350 reaktionerna 2
25351 reaktionära 1
25352 reaktionärerna 1
25353 reaktionärt 1
25354 reaktorer 8
25355 reaktorhaveri 1
25356 realinkomsten 1
25357 realism 1
25358 realismen 1
25359 realistisk 4
25360 realistiska 8
25361 realistiskt 10
25362 realitet 2
25363 realiteten 11
25364 realiteter 1
25365 realpolitiska 1
25366 realtid 1
25367 rebellerna 2
25368 recept 1
25369 reciprocal 1
25370 recirkulation 1
25371 recognised 1
25372 recovering 1
25373 recycling 1
25374 red 2
25375 reda 28
25376 redaktionella 2
25377 redan 503
25378 redare 1
25379 redares 1
25380 redarna 1
25381 redarnas 1
25382 redas 3
25383 rederi 1
25384 rederier 1
25385 rederiernas 1
25386 rederiet 2
25387 redigera 3
25388 redigerar 3
25389 redlighet 1
25390 redo 9
25391 redogjorde 2
25392 redogjort 4
25393 redogör 2
25394 redogöra 7
25395 redogörelse 5
25396 redogörelsen 1
25397 redogörelser 6
25398 redogörs 1
25399 redovisa 8
25400 redovisade 1
25401 redovisas 1
25402 redovisat 3
25403 redovisats 1
25404 redovisning 3
25405 redovisningskalkylerna 1
25406 redovisningsrubriker 1
25407 redovisningsskyldighet 1
25408 redskap 10
25409 reducera 4
25410 reducerar 1
25411 reduceras 6
25412 reducerat 3
25413 reducerats 1
25414 reducering 2
25415 reduceringen 1
25416 reell 8
25417 reella 8
25418 reellt 2
25419 referensbelopp 3
25420 referensbeloppen 1
25421 referensbibliotek 1
25422 referensen 5
25423 referenser 4
25424 referensfil 1
25425 referensfilen 2
25426 referenspunkt 3
25427 referensram 3
25428 referensramar 2
25429 referensramarna 2
25430 referera 1
25431 refererade 4
25432 refererar 3
25433 refereras 1
25434 reflektera 7
25435 reflektion 1
25436 reflektioner 1
25437 reflektionsarbete 3
25438 reflektionsarbeten 1
25439 reflektionslinje 1
25440 reflektionsplan 1
25441 reflex 1
25442 reflexion 1
25443 reflexionen 1
25444 reflexioner 1
25445 reform 60
25446 reform- 1
25447 reformansträngningar 1
25448 reformarbete 3
25449 reformarbetet 1
25450 reformatorn 1
25451 reformen 29
25452 reformens 6
25453 reformer 48
25454 reformera 14
25455 reformerade 1
25456 reformerar 3
25457 reformeras 6
25458 reformering 12
25459 reformeringen 11
25460 reformeringsmotor 1
25461 reformerna 19
25462 reformförfarande 1
25463 reformförslag 2
25464 reformförslagen 1
25465 reforminstrument 1
25466 reformister 1
25467 reformistisk 1
25468 reformistiska 11
25469 reformpaket 1
25470 reformprocess 4
25471 reformprocessen 7
25472 reformprogram 3
25473 reformprojektet 1
25474 reformsträvanden 1
25475 reformstämpel 1
25476 reformvilja 1
25477 reformvänlig 1
25478 reformvänliga 1
25479 reformåtgärder 1
25480 refuse 1
25481 regel 14
25482 regelbrott 1
25483 regelbunden 4
25484 regelbundenheten 1
25485 regelbundet 21
25486 regelbundna 6
25487 regellös 1
25488 regelmässig 1
25489 regelmässigt 2
25490 regeln 9
25491 regelrätt 1
25492 regelrätta 1
25493 regelsystem 1
25494 regelsystemet 1
25495 regelverk 22
25496 regelverken 1
25497 regelverket 9
25498 regera 1
25499 regerande 4
25500 regerandet 1
25501 regerar 1
25502 regerat 1
25503 regering 85
25504 regeringar 61
25505 regeringarna 41
25506 regeringarnas 7
25507 regeringars 2
25508 regeringen 120
25509 regeringens 20
25510 regerings 3
25511 regeringsbildning 1
25512 regeringsbildningen 9
25513 regeringschef 2
25514 regeringschefer 5
25515 regeringscheferna 9
25516 regeringschefernas 3
25517 regeringsfilosofin 1
25518 regeringsfunktioner 1
25519 regeringsföreträdare 1
25520 regeringsförfarande 1
25521 regeringsförhandlingarna 2
25522 regeringsförklaringen 1
25523 regeringskoalition 2
25524 regeringskoalitionens 1
25525 regeringskonferens 36
25526 regeringskonferensen 122
25527 regeringskonferensens 17
25528 regeringskonferenser 2
25529 regeringskritiker 1
25530 regeringslösningen 1
25531 regeringsmedlemmar 1
25532 regeringsmedlemmarna 1
25533 regeringsmedlemmars 1
25534 regeringsnivå 2
25535 regeringsorgan 1
25536 regeringsorganisationer 1
25537 regeringspartiet 4
25538 regeringsprogram 2
25539 regeringssamarbetets 1
25540 regeringssamarbetsnivå 1
25541 regeringsstrukturen 1
25542 regeringstjänstemän 1
25543 regeringsverksamheten 1
25544 regi 1
25545 regim 7
25546 regimen 8
25547 regimens 2
25548 regimer 4
25549 regimerna 1
25550 region 59
25551 regional 32
25552 regional- 1
25553 regionala 121
25554 regionalisering 1
25555 regionalister 1
25556 regionalplanering 1
25557 regionalplaneringspolitiken 1
25558 regionalpolitik 55
25559 regionalpolitiken 11
25560 regionalpolitikens 2
25561 regionalpolitiska 3
25562 regionalpresident 2
25563 regionalstöd 2
25564 regionalstödet 1
25565 regionalt 13
25566 regionen 72
25567 regionens 6
25568 regioner 145
25569 regionerna 83
25570 regionernas 10
25571 regioners 4
25572 regionnät 1
25573 register 10
25574 registrera 4
25575 registrerad 4
25576 registrerade 2
25577 registrerades 1
25578 registrerar 3
25579 registreras 3
25580 registrerat 1
25581 registrerats 1
25582 registrering 1
25583 registreringen 1
25584 registret 1
25585 regler 110
25586 reglera 14
25587 reglerad 2
25588 reglerade 6
25589 reglerande 3
25590 reglerandet 1
25591 reglerar 10
25592 regleras 13
25593 reglerat 2
25594 reglerats 2
25595 reglering 26
25596 regleringar 3
25597 regleringen 11
25598 regleringsförfarandet 1
25599 regleringskommitté 1
25600 reglerna 41
25601 reglernas 1
25602 regn 4
25603 regna 1
25604 regnade 1
25605 regnbågsringar 1
25606 regndroppsdiamanter 1
25607 regnet 2
25608 regnfloderna 1
25609 regnvatten 1
25610 regressiva 1
25611 reguljära 1
25612 rehabilitering 1
25613 rehabiliteringsprogram 1
25614 rejäl 1
25615 rejäla 3
25616 rejält 6
25617 reklam 6
25618 reklam- 1
25619 reklamdirektör 1
25620 reklamman 1
25621 reklamploj 1
25622 reklamvärldens 1
25623 rekognosceringsturer 1
25624 rekommendation 17
25625 rekommendationen 10
25626 rekommendationer 26
25627 rekommendationerna 19
25628 rekommendera 6
25629 rekommenderade 5
25630 rekommenderades 1
25631 rekommenderar 15
25632 rekommenderas 5
25633 rekommenderat 4
25634 rekonstruktion 2
25635 rekonstruktionsplan 1
25636 rekord 4
25637 rekordsnabb 1
25638 rekordtid 1
25639 rekreationslandskapet 1
25640 rekrytera 1
25641 rekryteringen 1
25642 rekryteringsmetoder 1
25643 rektor 1
25644 relaterade 3
25645 relateras 1
25646 relation 6
25647 relationen 1
25648 relationer 12
25649 relationerna 9
25650 relativ 6
25651 relativa 2
25652 relativisera 1
25653 relativt 18
25654 relevansen 1
25655 relevant 18
25656 relevanta 17
25657 reliable 1
25658 religion 7
25659 religionsanhängare 1
25660 religiös 2
25661 religiösa 3
25662 religiöst 2
25663 reliken 1
25664 reliker 2
25665 relikerna 1
25666 remiss 1
25667 remora 1
25668 remoran 1
25669 ren 27
25670 rena 24
25671 renar 1
25672 renare 6
25673 renas 1
25674 rengör 1
25675 rengöring 1
25676 rengöringen 1
25677 rengöringskrämer 1
25678 renhet 1
25679 rening 1
25680 reningsstationer 1
25681 reningsverk 2
25682 renligare 1
25683 renovera 1
25684 renoverar 1
25685 renovering 1
25686 renoveringen 1
25687 rensa 6
25688 rensar 1
25689 rensas 1
25690 rensat 2
25691 renskurat 1
25692 rensning 9
25693 rensningen 5
25694 rent 72
25695 rentav 8
25696 rentvättade 1
25697 renässans 1
25698 repade 1
25699 reparationerna 2
25700 reparera 6
25701 reparerat 1
25702 repet 1
25703 repknutar 1
25704 replikerna 1
25705 reportern 1
25706 representant 21
25707 representanten 15
25708 representantens 5
25709 representanter 4
25710 representanthuset 1
25711 representation 10
25712 representationen 2
25713 representationerna 1
25714 representativ 1
25715 representativa 6
25716 representativitet 3
25717 representativt 5
25718 representerade 3
25719 representerar 2
25720 representerat 1
25721 repression 1
25722 repressiva 1
25723 reproduktion 1
25724 reproduktionen 1
25725 reproduktiva 2
25726 reprulle 1
25727 republik 1
25728 republikanerna 4
25729 republikansk 1
25730 republikanska 1
25731 republiken 29
25732 republikens 6
25733 republikerna 2
25734 requis 2
25735 requérant 2
25736 resa 20
25737 resande 1
25738 resandet 1
25739 resans 1
25740 researrangörer 1
25741 researrangörernas 2
25742 resenärer 2
25743 reser 7
25744 reserv 3
25745 reservation 2
25746 reservationer 7
25747 reservationslöst 1
25748 reserven 1
25749 reserver 3
25750 reservera 1
25751 reserverad 1
25752 reserverade 4
25753 reserveras 1
25754 reserverats 1
25755 reservoarpenna 1
25756 reservoarpennor 1
25757 reservtrupper 1
25758 residens 1
25759 residuer 1
25760 resignera 1
25761 resklar 1
25762 resning 1
25763 resolut 2
25764 resolution 117
25765 resolutionen 81
25766 resolutionen.)Talmannen 1
25767 resolutionens 2
25768 resolutioner 26
25769 resolutionerna 6
25770 resolutionsförslag 36
25771 resolutionsförslagen 2
25772 resolutionsförslaget 14
25773 resolutionsförslagets 1
25774 resolutionstext 1
25775 resonanslåda 1
25776 resonemang 7
25777 resonemangen 2
25778 resonemanget 1
25779 resonera 1
25780 resonerade 2
25781 resonliga 1
25782 resor 4
25783 resource 1
25784 resp. 2
25785 respekt 78
25786 respektabel 1
25787 respektabelt 1
25788 respektabilitet 1
25789 respekten 34
25790 respektera 30
25791 respekterar 31
25792 respekteras 28
25793 respekterat 1
25794 respektfull 1
25795 respektingivande 2
25796 respektive 44
25797 respons 3
25798 responsibilise 1
25799 rest 5
25800 rest-Jugoslavien 1
25801 restaurang 2
25802 restaurangförbunden 1
25803 restaureringsarbetena 1
25804 reste 8
25805 resten 20
25806 rester 1
25807 resterande 4
25808 resterna 2
25809 restriktion 1
25810 restriktioner 2
25811 restriktionerna 3
25812 restriktiv 1
25813 restriktiva 1
25814 restriktivt 1
25815 rests 1
25816 restvara 1
25817 restämnen 1
25818 resultant 1
25819 resultat 146
25820 resultaten 37
25821 resultatet 42
25822 resultatinriktad 1
25823 resultatlista 1
25824 resultattavla 6
25825 resultattavlan 1
25826 resultatöversikt 4
25827 resultatöversikten 2
25828 resultera 1
25829 resulterade 3
25830 resulterar 8
25831 resulterat 4
25832 resurs 13
25833 resursbristen 1
25834 resursen 3
25835 resurser 114
25836 resurserna 36
25837 resursernas 2
25838 resursfrågor 1
25839 resursförbrukningskostnaderna 1
25840 resursfördelning 2
25841 resursförvaltning 1
25842 resurskrävande 1
25843 resursproblem 1
25844 resursslöseri 1
25845 resurstilldelning 1
25846 resväska 2
25847 resårer 1
25848 reta 1
25849 retar 1
25850 retirera 1
25851 retorik 12
25852 retroaktiv 1
25853 retroaktiva 3
25854 retroaktivitet 3
25855 retroaktiviteten 1
25856 retroaktivt 5
25857 retrospektiv 1
25858 reträtt 3
25859 returnerar 3
25860 rev 1
25861 revben 3
25862 revidera 8
25863 reviderade 3
25864 revideras 4
25865 revidering 17
25866 revideringar 1
25867 revideringen 10
25868 revideringsklausul 1
25869 revideringsklausulen 1
25870 revirstrider 1
25871 revision 6
25872 revisionen 1
25873 revisionsarbetskommittén 1
25874 revisionsarbetskommittés 1
25875 revisionsenheten 1
25876 revisionsfunktioner 1
25877 revisionsförklaring 1
25878 revisionsförklaringen 1
25879 revisionsroller 1
25880 revisionsrätten 13
25881 revisionsrättens 6
25882 revisionssystem 2
25883 revisionstjänst 2
25884 revisionstjänsten 2
25885 revisionsuppföljning 1
25886 revolution 6
25887 revolutionen 3
25888 revolutioner 1
25889 revolutionslandet 1
25890 revolutionsregeringens 1
25891 revolutionär 3
25892 revolutionära 2
25893 revolver 1
25894 ribban 1
25895 rida 2
25896 riddare 3
25897 ridå 1
25898 ridån 1
25899 riggade 1
25900 rights 1
25901 rigiditeten 1
25902 rigorös 1
25903 rigorösa 3
25904 rigoröst 4
25905 rik 3
25906 rika 19
25907 rikare 3
25908 rikaste 5
25909 rikedom 7
25910 rikedomar 7
25911 rikedomarna 3
25912 rikedomen 6
25913 riket 2
25914 riklig 5
25915 rikligt 1
25916 riksdagen 1
25917 riksdagens 1
25918 riksdagsledamöter 1
25919 rikt 4
25920 rikta 26
25921 riktad 4
25922 riktade 15
25923 riktades 1
25924 riktar 12
25925 riktas 10
25926 riktat 3
25927 riktats 2
25928 riktig 23
25929 riktiga 7
25930 riktige 1
25931 riktigt 79
25932 riktlinje 2
25933 riktlinjen 2
25934 riktlinjer 85
25935 riktlinjerna 42
25936 riktlinjernas 3
25937 riktning 59
25938 riktningar 1
25939 riktningarna 2
25940 riktningen 15
25941 riktpunkter 2
25942 rimlig 11
25943 rimliga 14
25944 rimligare 1
25945 rimligen 2
25946 rimligt 16
25947 rimligtvis 1
25948 rimmar 1
25949 ring 2
25950 ringa 11
25951 ringakta 1
25952 ringde 8
25953 ringen 1
25954 ringer 6
25955 ringklockan 1
25956 ringlade 1
25957 ringt 1
25958 rinner 1
25959 ris 2
25960 risk 34
25961 riskabel 3
25962 riskanalys 3
25963 riskavfall 1
25964 riskbedömning 3
25965 riskbedömningen 1
25966 risken 39
25967 risker 32
25968 riskera 7
25969 riskerade 1
25970 riskerar 42
25971 riskerna 17
25972 riskexponering 1
25973 riskfaktor 1
25974 riskfritt 1
25975 riskfylld 2
25976 riskfyllda 4
25977 riskfyllt 2
25978 riskförebyggande 2
25979 riskhantering 5
25980 riskhanteringsfunktion 1
25981 riskkapital 6
25982 riskkommunikation 2
25983 risknivå 1
25984 riskspridning 1
25985 riskspridningsprincipen 1
25986 riskspridningsregler 2
25987 risktagande 2
25988 risktagarna 1
25989 riskuppgifterna 1
25990 riskutvecklingen 1
25991 riskvilligt 1
25992 riskvärdering 3
25993 riskzonen 2
25994 riste 1
25995 ritat 1
25996 ritualbärare 1
25997 rituell 1
25998 rituella 1
25999 riva 1
26000 rivalen 1
26001 rivs 1
26002 ro 7
26003 roade 4
26004 roar 2
26005 roat 2
26006 robusta 1
26007 rocken 1
26008 rockfickan 1
26009 rockskört 1
26010 roder 1
26011 rodret 1
26012 roffa 1
26013 rofylld 1
26014 roliga 1
26015 roligt 12
26016 roll 221
26017 rollen 12
26018 roller 4
26019 roman 1
26020 romantiken 1
26021 romantiska 1
26022 romarna 2
26023 romarnas 1
26024 romer 6
26025 romerbefolkningen 1
26026 romergruppen 1
26027 romerna 2
26028 romernas 1
26029 ropa 2
26030 ropade 6
26031 ropande 1
26032 ropar 4
26033 ropet 2
26034 ros 3
26035 rosa 1
26036 rosafärgad 1
26037 rosenröd 1
26038 rosenrött 1
26039 rosig 1
26040 rosor 1
26041 rosorna 2
26042 rostade 3
26043 rostar 1
26044 rostat 1
26045 rostbildning 1
26046 rostig 2
26047 rostiga 1
26048 rota 1
26049 rotade 1
26050 rotat 1
26051 rotation 1
26052 rotelement 1
26053 rotelementet 1
26054 roten 1
26055 rotsystem 1
26056 rott 1
26057 round 1
26058 rovfiske 1
26059 rubba 1
26060 rubbar 1
26061 rubbas 1
26062 rubbat 1
26063 rubbats 1
26064 rubbningarna 1
26065 rubrik 14
26066 rubriken 3
26067 rubriker 2
26068 rubrikerna 1
26069 ruelse 1
26070 ruffig 1
26071 ruffiga 1
26072 rufsigt 1
26073 rugbybrede 1
26074 ruin 2
26075 ruiner 2
26076 ruinerad 1
26077 ruineras 1
26078 ruinerna 1
26079 ruljangsen 1
26080 rullade 2
26081 rullande 1
26082 rullar 4
26083 rullat 2
26084 rullats 1
26085 rullstol 1
26086 rullstolen 1
26087 rullstolsburna 1
26088 rum 135
26089 rumlade 1
26090 rummel 1
26091 rummet 16
26092 rumänsk 1
26093 rumänska 4
26094 rund 1
26095 runda 8
26096 rundabordskonferens 1
26097 rundan 3
26098 rundor 2
26099 rundresa 3
26100 rundresan 1
26101 rundtur 1
26102 runt 45
26103 runtom 2
26104 rusa 3
26105 rusade 11
26106 rusande 1
26107 rusar 4
26108 ruskig 1
26109 rusta 2
26110 rustad 2
26111 rustningsproblemets 1
26112 rutan 1
26113 rutig 1
26114 rutin 2
26115 rutinen 2
26116 rutiner 12
26117 rutinerna 3
26118 rutinmässiga 2
26119 rutmönster 1
26120 rutnät 1
26121 rutnätets 2
26122 ruttna 3
26123 ruttnade 1
26124 ruttnande 1
26125 ruvade 3
26126 ruvande 2
26127 ryck 1
26128 rycka 2
26129 rycker 1
26130 ryckig 1
26131 ryckigt 1
26132 ryckte 3
26133 ryckts 1
26134 rygg 6
26135 rygga 2
26136 ryggar 1
26137 ryggen 10
26138 ryggmusklerna 1
26139 ryggrad 2
26140 ryggraden 1
26141 ryktas 1
26142 ryktbarhet 1
26143 rykte 7
26144 rykten 2
26145 ryktena 1
26146 rymde 2
26147 rymden 7
26148 rymdmonster 1
26149 rymdåldern 1
26150 rymma 2
26151 rymmer 2
26152 ryms 1
26153 rynkor 1
26154 rysk 1
26155 ryska 15
26156 ryske 9
26157 rysning 1
26158 ryssar 1
26159 ryssarna 1
26160 rytm 3
26161 rytmiskt 1
26162 räcka 16
26163 räcker 59
26164 räckhåll 2
26165 räcks 1
26166 räckte 13
26167 räckvidd 6
26168 rädd 13
26169 rädda 30
26170 räddade 2
26171 räddades 1
26172 räddande 1
26173 räddar 2
26174 räddas 1
26175 räddat 1
26176 räddats 1
26177 räddning 3
26178 räddningen 2
26179 räddningshelikoptrar 2
26180 räddningsnivåer 1
26181 räddningstjänst 1
26182 räddningstjänster 1
26183 rädsla 10
26184 rädslan 5
26185 räkenskap 2
26186 räkenskaper 1
26187 räkenskaperna 7
26188 räkenskapsansvariga 1
26189 räkenskapssystemet 1
26190 räkenskapsår 1
26191 räkna 25
26192 räknade 2
26193 räknar 39
26194 räknas 7
26195 räknat 8
26196 räknats 1
26197 räkneexempel 1
26198 räkning 31
26199 räkningar 1
26200 räkningen 2
26201 räls 1
26202 räntan 1
26203 räntehöjning 1
26204 ränteintäkter 1
26205 ränteutgifter 1
26206 räntor 1
26207 räntorna 1
26208 rät 1
26209 räta 1
26210 rätas 1
26211 rätt 282
26212 rätta 73
26213 rättade 1
26214 rättades 1
26215 rättan 1
26216 rättar 1
26217 rättas 3
26218 rättats 2
26219 rättegång 6
26220 rättegångar 2
26221 rättegången 1
26222 rättegångsprocesser 1
26223 rätteligen 2
26224 rättelse 1
26225 rätten 72
26226 rättens 1
26227 rättfram 2
26228 rättframt 2
26229 rättfärdiga 5
26230 rättfärdigande 1
26231 rättfärdiganden 1
26232 rättfärdigandet 1
26233 rättfärdigar 4
26234 rättfärdigas 2
26235 rättfärdigat 1
26236 rättfärdigt 1
26237 rättighet 23
26238 rättigheten 1
26239 rättigheter 276
26240 rättigheterna 174
26241 rättigheternas 5
26242 rättigheters 1
26243 rättighetsinnehavarna 2
26244 rättighetsstadgor 1
26245 rättmätig 2
26246 rättmätiga 2
26247 rättmätigt 2
26248 rättrogna 1
26249 rättrådigheten 1
26250 rätts- 1
26251 rättsakt 4
26252 rättsakter 3
26253 rättsdefinition 1
26254 rättsförluster 1
26255 rättshjälp 20
26256 rättshjälpen 4
26257 rättsinniga 1
26258 rättsinstanser 2
26259 rättsinstanserna 1
26260 rättskaffens 2
26261 rättskipning 7
26262 rättskipningssystemet 1
26263 rättskultur 1
26264 rättskulturen 1
26265 rättslig 55
26266 rättsliga 164
26267 rättsligt 36
26268 rättsläget 3
26269 rättsområde 2
26270 rättsordning 1
26271 rättsordningen 2
26272 rättsosäkerhet 2
26273 rättspraxis 3
26274 rättsprincip 1
26275 rättsprinciper 1
26276 rättsprocess 1
26277 rättsprocessen 2
26278 rättsregler 1
26279 rättsreglerna 1
26280 rättssamarbetet 1
26281 rättssekreterare 1
26282 rättsskipande 3
26283 rättsskipning 2
26284 rättsskipningen 2
26285 rättsskydd 1
26286 rättsskyddsområdet 1
26287 rättsstat 5
26288 rättsstaten 4
26289 rättsstatens 2
26290 rättsstatliga 1
26291 rättsstatlighet 2
26292 rättsstatsprincip 1
26293 rättsstatsprincipen 2
26294 rättsstatus 1
26295 rättsstödet 1
26296 rättssystem 17
26297 rättssystemen 8
26298 rättssystemet 7
26299 rättssäkerhet 15
26300 rättssäkerheten 8
26301 rättstillämpningen 1
26302 rättstjänst 1
26303 rättstjänsten 1
26304 rättstraditionen 1
26305 rättstraditioner 2
26306 rättsuppfattningen 1
26307 rättsutskottet 1
26308 rättsutskottets 1
26309 rättsväsen 1
26310 rättsväsende 4
26311 rättsväsendet 3
26312 rätttsliga 1
26313 rättvis 28
26314 rättvisa 85
26315 rättvisan 10
26316 rättvisans 2
26317 rättvisare 2
26318 rättvisebehov 1
26319 rättvisefrågor 1
26320 rättvisekriterier 1
26321 rättvist 29
26322 rättänkande 1
26323 rå 1
26324 råa 1
26325 råare 1
26326 råd 38
26327 råda 22
26328 rådande 8
26329 rådde 8
26330 rådens 2
26331 råder 71
26332 rådet 504
26333 rådets 268
26334 rådfråga 3
26335 rådfrågades 2
26336 rådfrågar 2
26337 rådfrågat 2
26338 rådfrågats 2
26339 rådfrågningar 1
26340 rådfrågningsprocessen 1
26341 rådgivande 14
26342 rådgivare 5
26343 rådgivarna 1
26344 rådgivarnas 1
26345 rådgivning 7
26346 rådgivningen 1
26347 rådgivningsnätverk 1
26348 rådgivningsverksamhet 1
26349 rådgör 1
26350 rådighet 1
26351 råds 2
26352 rådsbeslut 1
26353 rådsbeslutet 1
26354 rådsförsamlingar 1
26355 rådsgruppen 1
26356 rådslag 3
26357 rådsledamöterna 1
26358 rådsmedlemmar 1
26359 rådsministrar 1
26360 rådsmötena 1
26361 rådsmötet 9
26362 rådsordförande 55
26363 rådsordföranden 18
26364 rådsordförandens 3
26365 rådsordförandeskapet 3
26366 rådsordförandeskapets 1
26367 rådsrepresentanternas 1
26368 rådsresolution 1
26369 rådstoppmötet 1
26370 rågata 1
26371 råkade 5
26372 råkar 3
26373 råkat 2
26374 råmaterial 3
26375 råmärken 1
26376 rånares 1
26377 rånkupp 1
26378 råolja 3
26379 råskinn 1
26380 rått 4
26381 råttan 1
26382 råttor 1
26383 råvara 1
26384 råvaror 1
26385 råvarorna 1
26386 råvaruproducenter 1
26387 référendaire 1
26388 röd 8
26389 röda 19
26390 rödgröna 1
26391 rödhårig 1
26392 rödklädda 1
26393 rödrutig 1
26394 rödvin 1
26395 rödögda 1
26396 rök 2
26397 röka 1
26398 röken 1
26399 röker 2
26400 rökgrå 1
26401 rökmoln 1
26402 rökningen 1
26403 rökpuffar 1
26404 rökridåer 1
26405 rökte 5
26406 rönt 1
26407 rönte 1
26408 rör 113
26409 röra 16
26410 röran 1
26411 rörande 64
26412 röras 1
26413 rörde 11
26414 rörelse 11
26415 rörelsehindrade 1
26416 rörelsen 3
26417 rörelser 8
26418 rörelserna 1
26419 rören 1
26420 rörig 1
26421 rörigt 3
26422 rörlig 2
26423 rörliga 3
26424 rörlighet 30
26425 rörligheten 18
26426 rört 4
26427 röst 42
26428 rösta 112
26429 röstade 37
26430 röstades 3
26431 röstar 36
26432 röstas 4
26433 röstat 40
26434 röstats 1
26435 rösten 6
26436 röster 18
26437 rösterna 2
26438 röstförklaring 7
26439 röstförklaringar 1
26440 röstförklaringarna 1
26441 röstkapacitet 1
26442 röstlista 1
26443 röstresultat 1
26444 rösträtt 4
26445 rösträtten 3
26446 röstsystem 2
26447 röstsystemet 2
26448 röstsystemsfråga 1
26449 röstviktning 3
26450 rött 7
26451 rötter 5
26452 rötterna 2
26453 rövats 1
26454 s 3
26455 s'il 1
26456 s. 1
26457 s.16 1
26458 s.k. 16
26459 sa 94
26460 sabeltandad 1
26461 sade 249
26462 sades 3
26463 safety-protokollet 1
26464 sagan 1
26465 sagda 1
26466 sagt 159
26467 sagts 31
26468 sak 114
26469 sak- 3
26470 saken 36
26471 sakens 4
26472 saker 106
26473 sakerna 7
26474 sakernas 2
26475 sakfrågan 3
26476 sakfrågor 2
26477 sakförhållanden 1
26478 sakförhållandena 1
26479 sakinnehållet 1
26480 sakkunnig 1
26481 sakkunniga 6
26482 sakkunskap 4
26483 sakkunskapen 1
26484 sakkännedom 2
26485 saklig 1
26486 sakliga 2
26487 sakligt 1
26488 sakna 1
26489 saknade 8
26490 saknaden 1
26491 saknades 3
26492 saknar 34
26493 saknas 58
26494 saknat 2
26495 saknats 1
26496 sakområden 1
26497 sakområdet 1
26498 sakproblem 1
26499 sakta 14
26500 sakupplysning 1
26501 sal 1
26502 salen 2
26503 salinarbetare 1
26504 salladsblad 1
26505 saltdofter 1
26506 saltvatten 1
26507 salu 2
26508 saluföra 2
26509 saluförande 1
26510 saluförandet 1
26511 saluförde 1
26512 saluföringen 3
26513 saluföringsfrågorna 1
26514 saluföringskostnaderna 1
26515 saluförs 2
26516 samarbeta 27
26517 samarbetar 12
26518 samarbetat 3
26519 samarbete 168
26520 samarbetet 86
26521 samarbetets 3
26522 samarbets- 3
26523 samarbetsanda 4
26524 samarbetsavtal 4
26525 samarbetsavtalet 3
26526 samarbetsbetonat 1
26527 samarbetskapacitet 1
26528 samarbetsklimat 1
26529 samarbetskommittén 1
26530 samarbetsländerna 1
26531 samarbetsmodell 1
26532 samarbetsområden 1
26533 samarbetsområdena 2
26534 samarbetsorganisation 1
26535 samarbetspartner 1
26536 samarbetspolitik 5
26537 samarbetspolitiken 5
26538 samarbetsprincipen 1
26539 samarbetsprocess 1
26540 samarbetsprogram 1
26541 samarbetsprojekt 3
26542 samarbetsprojekten 1
26543 samarbetsramen 1
26544 samarbetsstrategi 1
26545 samarbetssätt 1
26546 samarbetsutveckling 1
26547 samarbetsvilja 1
26548 samarbetsvilliga 1
26549 samband 138
26550 sambanden 2
26551 sambandet 4
26552 samexistens 7
26553 samexistensen 1
26554 samfinansierades 1
26555 samfinansieras 1
26556 samfinansiering 2
26557 samfinansieringen 1
26558 samfund 1
26559 samfunden 2
26560 samfundet 11
26561 samfundets 3
26562 samförstånd 21
26563 samförståndspolitik 1
26564 samhälle 50
26565 samhällelig 2
26566 samhälleliga 3
26567 samhällen 33
26568 samhällena 5
26569 samhälles 4
26570 samhället 79
26571 samhällets 15
26572 samhällsaktörer 1
26573 samhällsansvar 1
26574 samhällsekonomin 1
26575 samhällsekonomisk 1
26576 samhällsekonomiska 3
26577 samhällsfaktor 1
26578 samhällsfientliga 1
26579 samhällsgrupperna 1
26580 samhällsklasser 1
26581 samhällskostnaderna 1
26582 samhällsliv 2
26583 samhällslivet 1
26584 samhällsmedborgare 1
26585 samhällsmodell 1
26586 samhällsmodellen 3
26587 samhällsomfattande 11
26588 samhällsomgivningen 1
26589 samhällsområden 1
26590 samhällspolitiska 1
26591 samhällsservicen 1
26592 samhällsstöd 1
26593 samhällssystem 1
26594 samhällsteori 1
26595 samhällsvärde 1
26596 samhörande 1
26597 samhörigheten 1
26598 samklang 2
26599 samla 22
26600 samlad 2
26601 samlade 13
26602 samlades 3
26603 samlar 3
26604 samlarfordon 1
26605 samlarmani 1
26606 samlas 6
26607 samlat 9
26608 samlats 5
26609 samlevnad 3
26610 samlevnaden 1
26611 samlevnadsformer 1
26612 samling 7
26613 samlingsplatser 1
26614 samma 289
26615 sammalunda 1
26616 samman 56
26617 sammanbindande 1
26618 sammanblanda 1
26619 sammanblandning 2
26620 sammanboende 1
26621 sammanbrott 1
26622 sammanbunden 1
26623 sammandrabbning 1
26624 sammandrag 1
26625 sammanfalla 1
26626 sammanfallande 1
26627 sammanfallanden 1
26628 sammanfaller 5
26629 sammanfatta 8
26630 sammanfattade 1
26631 sammanfattande 1
26632 sammanfattar 4
26633 sammanfattas 3
26634 sammanfattat 2
26635 sammanfattning 10
26636 sammanfattningar 1
26637 sammanfattningen 1
26638 sammanfattningsvis 6
26639 sammanflätade 2
26640 sammanfogas 1
26641 sammanfogat 1
26642 sammanför 1
26643 sammanföra 5
26644 sammanföras 1
26645 sammanförde 1
26646 sammanhang 85
26647 sammanhangen 2
26648 sammanhanget 49
26649 sammanhopningen 2
26650 sammanhängande 10
26651 sammanhänger 1
26652 sammanhållande 2
26653 sammanhållen 2
26654 sammanhållning 63
26655 sammanhållningen 45
26656 sammanhållningsfonden 1
26657 sammanhållningsländerna 2
26658 sammanhållningspolitik 3
26659 sammanhållningspolitiken 2
26660 sammanhållningspolitikens 2
26661 sammanhållningsprocessen 2
26662 sammanhörande 2
26663 sammanjämka 2
26664 sammanjämkar 1
26665 sammankalla 5
26666 sammankallande 2
26667 sammankallandet 4
26668 sammankallas 1
26669 sammankomst 1
26670 sammankomster 1
26671 sammankomsterna 1
26672 sammankoppla 1
26673 sammankopplade 2
26674 sammanlagd 1
26675 sammanlagda 3
26676 sammanlagt 4
26677 sammanlänka 1
26678 sammanlänkade 1
26679 sammansatt 7
26680 sammanslaget 1
26681 sammanslagning 3
26682 sammanslagningar 6
26683 sammanslagningen 4
26684 sammanslagningsvåg 1
26685 sammanslutning 2
26686 sammanslutningar 6
26687 sammanslutningarna 2
26688 sammanslutnings 1
26689 sammansmältningens 1
26690 sammanställa 2
26691 sammanställd 1
26692 sammanställde 1
26693 sammanställer 1
26694 sammanställning 6
26695 sammanställningen 4
26696 sammanställs 1
26697 sammanställt 2
26698 sammanställts 1
26699 sammansvärjning 1
26700 sammansättning 6
26701 sammansättningen 6
26702 sammanträda 3
26703 sammanträdde 1
26704 sammanträde 30
26705 sammanträden 4
26706 sammanträdena 4
26707 sammanträder 4
26708 sammanträdesperiod 7
26709 sammanträdesperioden 2
26710 sammanträdesperiodens 1
26711 sammanträdesperioder 1
26712 sammanträdesperioderna 1
26713 sammanträdesrum 1
26714 sammanträdessessionen 1
26715 sammanträdestakten 1
26716 sammanträdet 25
26717 sammanträdets 1
26718 sammanträffande 1
26719 sammanträffanden 1
26720 sammanträtt 1
26721 sammetsdraperade 1
26722 sammetsstol 1
26723 samordna 26
26724 samordnad 11
26725 samordnade 13
26726 samordnande 2
26727 samordnar 2
26728 samordnare 4
26729 samordnarna 1
26730 samordnas 5
26731 samordnat 3
26732 samordnats 1
26733 samordning 60
26734 samordningen 25
26735 samordningsaspekt 1
26736 samordningsförfarandet 1
26737 samordningsförmåga 1
26738 samordningsmekanismer 1
26739 samordningsmetod 1
26740 samordningsproblem 1
26741 samordningsprocess 1
26742 samordningsstruktur 1
26743 samriskföretag 2
26744 samråd 19
26745 samråda 3
26746 samråden 2
26747 samrådet 2
26748 samrådsakt 1
26749 samrådsarbete 1
26750 samrådsdirektiv 1
26751 samrådsdokumentet 1
26752 samrådsforum 1
26753 samrådsförfarande 1
26754 samrådsförfaranden 1
26755 samrådsförfarandet 1
26756 samrådsförslaget 1
26757 samrådskommittéer 1
26758 samrådsprocess 1
26759 samrådsprocessen 1
26760 samrådsrättigheter 1
26761 samsats 1
26762 samspel 1
26763 samspelet 2
26764 samspråk 1
26765 samstämmig 6
26766 samstämmiga 3
26767 samstämmighet 63
26768 samstämmigheten 21
26769 samstämmighetsobservatorium 1
26770 samstämmighetspolitiken 1
26771 samstämmighetsprocessen 1
26772 samstämmighetsövervakning 1
26773 samstämmigt 7
26774 samstämt 1
26775 samsyn 5
26776 samt 228
26777 samtal 27
26778 samtala 2
26779 samtalar 1
26780 samtalen 12
26781 samtalet 5
26782 samtalspartner 3
26783 samtalsrundan 1
26784 samtalssvårigheter 1
26785 samtalsämne 1
26786 samtida 1
26787 samtidens 1
26788 samtidighet 1
26789 samtidigt 188
26790 samtliga 91
26791 samtycke 17
26792 samtycker 3
26793 samtyckesförfarandet 2
26794 samtyckt 1
26795 samvarotid 1
26796 samverka 6
26797 samverkan 5
26798 samverkande 1
26799 samverkar 2
26800 samvete 1
26801 samveten 3
26802 samvetet 3
26803 samvetsgranna 1
26804 samvetslös 1
26805 samvetsskäl 1
26806 sandaler 1
26807 sanden 1
26808 sandtag 1
26809 sanera 4
26810 sanerats 1
26811 saneringen 8
26812 saneringsarbete 1
26813 sanitär 2
26814 sanitära 3
26815 sanka 1
26816 sanktion 1
26817 sanktionen 1
26818 sanktioner 29
26819 sanktionera 2
26820 sanktionerad 1
26821 sanktionerna 7
26822 sanktionspolitik 1
26823 sanktionssystem 2
26824 sanktionssystemet 1
26825 sann 2
26826 sanna 1
26827 sannerligen 12
26828 sanning 4
26829 sanningen 13
26830 sanningens 1
26831 sannings- 1
26832 sannolika 1
26833 sannolikhet 5
26834 sannolikheten 1
26835 sannolikhetskalkyl 1
26836 sannolikt 15
26837 sansad 1
26838 sansat 2
26839 sant 45
26840 sargande 1
26841 sarkastisk 1
26842 satellit 2
26843 satelliter 1
26844 satellitteve 1
26845 satellitövervakning 2
26846 satsa 24
26847 satsade 1
26848 satsar 6
26849 satsas 3
26850 satsat 3
26851 satsats 1
26852 satsning 8
26853 satsningar 4
26854 satsningen 3
26855 satt 52
26856 satta 3
26857 satte 24
26858 sattes 4
26859 satts 6
26860 scale 1
26861 scen 1
26862 scenarbetare 1
26863 scenarier 3
26864 scenario 2
26865 scenarior 1
26866 scenariot 2
26867 scenen 4
26868 scener 1
26869 schablonmässigt 1
26870 schackbräde 1
26871 schema 3
26872 schemat 3
26873 schizofren 1
26874 schweiziska 2
26875 scientifiques 1
26876 scones 1
26877 sconesen 1
26878 scoreboard 1
26879 se 512
26880 securities 2
26881 sedan 344
26882 sedda 1
26883 seder 1
26884 sedlar 2
26885 sedlarna 2
26886 sedligt 1
26887 sedvanliga 3
26888 sedvanor 1
26889 seg 2
26890 segdraget 1
26891 segel 1
26892 segelbara 1
26893 segelfartyg 1
26894 segelleden 1
26895 seger 7
26896 segern 3
26897 segla 5
26898 seglade 4
26899 seglar 14
26900 seglat 1
26901 seglen 1
26902 seglingen 1
26903 segment 1
26904 segra 1
26905 segrat 1
26906 seismisk 1
26907 seismiska 1
26908 sekel 11
26909 sekellång 1
26910 sekellöst 1
26911 sekelskifte 1
26912 sekelskiftet 1
26913 sekelslutet 1
26914 sekler 1
26915 seklerna 1
26916 seklers 1
26917 seklet 2
26918 sekretariat 4
26919 sekretariatet 1
26920 sekreterare 3
26921 sekretess 6
26922 sekretessbelagd 1
26923 sekretessbelagda 3
26924 sekretessbelägga 1
26925 sekretessbelägger 1
26926 sekretessen 1
26927 sekretesshänsynen 1
26928 sektion 3
26929 sektor 39
26930 sektorer 46
26931 sektorerna 11
26932 sektoriell 3
26933 sektoriella 2
26934 sektorinriktad 2
26935 sektorinriktade 1
26936 sektorintressen 1
26937 sektorn 43
26938 sektorns 10
26939 sektorpolitik 1
26940 sektors 1
26941 sektorsanalys 1
26942 sektorsfråga 1
26943 sektorsinriktat 1
26944 sektorsspecifika 1
26945 sektorsövergripande 2
26946 sekulariserade 1
26947 sekund 4
26948 sekunder 5
26949 sekundärprocesser 1
26950 sekundärrätten 1
26951 sekundärtransvestit 1
26952 seldon 1
26953 selektiv 5
26954 selektiva 6
26955 selektivitet 1
26956 selektivt 8
26957 semantisk 1
26958 semester 7
26959 semesterfirare 1
26960 semesterfirarna 1
26961 semestertider 1
26962 semestra 1
26963 semestrar 1
26964 semestrarna 1
26965 seminarier 1
26966 seminarierna 1
26967 seminariet 1
26968 seminarium 3
26969 sen 18
26970 sena 3
26971 senare 104
26972 senareläggas 2
26973 senareläggning 1
26974 senast 19
26975 senaste 173
26976 senat 2
26977 senaten 2
26978 senator 4
26979 senatorer 1
26980 senfärdig 1
26981 sensibilitet 1
26982 sent 30
26983 sentimentalitet 1
26984 separat 5
26985 separata 7
26986 separatism 1
26987 separerade 1
26988 september 27
26989 ser 255
26990 sera 1
26991 serb 1
26992 serber 16
26993 serberna 4
26994 serbisk 1
26995 serbiska 7
26996 serie 8
26997 seriefält 1
26998 seriesläppområde 1
26999 seriös 5
27000 seriösa 6
27001 seriösare 1
27002 seriöst 20
27003 servats 1
27004 servera 3
27005 serverades 1
27006 serverar 1
27007 serveringsfat 1
27008 service 30
27009 serviceföretag 1
27010 servicekort 1
27011 servicekvalitet 2
27012 servicen 15
27013 servicenivå 1
27014 servicens 1
27015 servicenätverk 1
27016 ses 32
27017 session 20
27018 sessionen 20
27019 sessioner 3
27020 sessionerna 1
27021 sessionstiden 1
27022 sessionstjänsten 1
27023 sett 134
27024 setts 1
27025 sex 48
27026 sex- 1
27027 sexismen 1
27028 sexmånadersperiod 3
27029 sextio 2
27030 sextiotalet 4
27031 sextiotusenmannastyrkan 1
27032 sextiotvå 1
27033 sexton 4
27034 sextumskanonerna 2
27035 sexturismen 1
27036 sexuell 2
27037 sexuella 3
27038 sexuellt 2
27039 sexvärt 1
27040 sexårsdag 1
27041 sexårsperiod 1
27042 sfär 2
27043 sfärer 1
27044 shall 1
27045 sharing 1
27046 sherry 1
27047 shilling 1
27048 shipping 1
27049 shorts 2
27050 shownummer 1
27051 si 1
27052 sicilianska 1
27053 sida 141
27054 sidan 195
27055 sidans 1
27056 siden 1
27057 sidenklänning 1
27058 sidenträ 1
27059 sidfilnamn.bak.htm 1
27060 sidfot 1
27061 sidfotsektion 1
27062 sidhuvud 1
27063 sidhuvudsektion 1
27064 sidoblick 1
27065 sidoeffekter 1
27066 sidor 27
27067 sidorna 7
27068 siffermässiga 1
27069 siffra 7
27070 siffran 1
27071 siffror 19
27072 siffrorna 13
27073 sig 1694
27074 signal 19
27075 signalen 2
27076 signaler 7
27077 signalerar 2
27078 signerade 1
27079 signerar 1
27080 signerat 1
27081 signifikant 1
27082 signifikativt 1
27083 signum 1
27084 sikt 62
27085 sikta 2
27086 siktade 1
27087 siktar 6
27088 sikte 7
27089 siktet 1
27090 sill 1
27091 sillhuvuden 2
27092 silver 2
27093 silver- 1
27094 silvergarnityr 1
27095 silverglänsande 1
27096 silverräv 1
27097 silversiklar 1
27098 silverskimrande 1
27099 silvertråden 1
27100 simma 1
27101 simpel 2
27102 simpla 1
27103 simulatorer 2
27104 sin 597
27105 sina 433
27106 sinad 1
27107 sine 5
27108 singel 1
27109 sinnade 1
27110 sinnat 1
27111 sinne 2
27112 sinnelag 3
27113 sinnen 3
27114 sinnena 1
27115 sinnesrörelse 2
27116 sinnesstämning 1
27117 sinom 2
27118 sinsemellan 9
27119 sir 3
27120 sist 46
27121 sista 103
27122 siste 2
27123 sistnämnda 11
27124 sistnämndas 1
27125 sitt 347
27126 sitta 15
27127 sittande 1
27128 sittbad 1
27129 sitter 31
27130 sittning 2
27131 situation 127
27132 situationen 176
27133 situationens 6
27134 situationer 30
27135 situationerna 1
27136 sjabblar 1
27137 sjok 1
27138 sju 26
27139 sjudande 1
27140 sjuhundra 2
27141 sjuk 10
27142 sjuk- 2
27143 sjuka 3
27144 sjukdom 10
27145 sjukdomar 12
27146 sjukdomen 8
27147 sjukdomens 2
27148 sjukdomsbekämpning 1
27149 sjukdomsskydd 1
27150 sjukförsäkring 1
27151 sjukhus 9
27152 sjukhusen 1
27153 sjukhuset 7
27154 sjukhusplatserna 1
27155 sjukligt 2
27156 sjukvård 3
27157 sjukvården 1
27158 sjukvårdens 1
27159 sjukvårds- 1
27160 sjukvårdsanläggningar 1
27161 sjukvårdsbudgeten 1
27162 sjukvårdsfrågorna 1
27163 sjukvårdspolitik 1
27164 sjunde 5
27165 sjunga 1
27166 sjungande 1
27167 sjunger 1
27168 sjunka 9
27169 sjunkande 1
27170 sjunker 3
27171 sjunkit 9
27172 sjunkna 4
27173 sjutton 2
27174 sjuttonde 1
27175 sjuårsperiod 2
27176 själ 7
27177 själar 2
27178 själen 2
27179 själlösa 1
27180 själv 204
27181 själva 240
27182 självaktning 1
27183 självaste 1
27184 självbedrägeri 1
27185 självbedrägerier 1
27186 självbelåtenhet 1
27187 självbelåtne 1
27188 självbestämmande 6
27189 självbiografi 3
27190 självbärande 2
27191 självfallet 7
27192 självförnöjelse 1
27193 självförsörjande 2
27194 självförtroendet 1
27195 självförvaltande 1
27196 självförvållade 1
27197 självhjälp 3
27198 självklar 7
27199 självklara 4
27200 självklarhet 6
27201 självklart 49
27202 självkostnadspriser 1
27203 självkänsla 1
27204 självlysande 1
27205 självmant 1
27206 självmedlidande 1
27207 självmord 1
27208 självplågeri 1
27209 självrespekt 1
27210 självstympning 1
27211 självstyrande 6
27212 självstyre 2
27213 självstyrelse 3
27214 självstyrelsens 1
27215 självstyrelseorganen 1
27216 självstyret 1
27217 självständig 6
27218 självständiga 8
27219 självständighet 5
27220 självständigheten 1
27221 självständighetsdagen 1
27222 självständighetsfesten 1
27223 självständighetsfirandet 1
27224 självständighetsprocess 1
27225 självständighetsrörelsen 1
27226 självständigt 10
27227 självsäkert 3
27228 självt 22
27229 självtillit 1
27230 självtäkt 1
27231 självverkande 1
27232 självändamål 4
27233 sjätte 21
27234 sjättedel 1
27235 sjöar 3
27236 sjöarna 1
27237 sjöcertifikat 1
27238 sjöd 1
27239 sjödugligt 1
27240 sjöfarandes 1
27241 sjöfarten 1
27242 sjöfartens 1
27243 sjöfartsinspektionen 1
27244 sjöfartsmyndigheter 1
27245 sjöfartsområdena 1
27246 sjöfartsorganisationen 2
27247 sjöfartssektorn 3
27248 sjöfolk 1
27249 sjögående 1
27250 sjöman 5
27251 sjömannamässigt 1
27252 sjömannen 1
27253 sjömän 3
27254 sjömännen 3
27255 sjön 11
27256 sjöng 3
27257 sjönk 10
27258 sjöovärdiga 1
27259 sjörätt 1
27260 sjöss 7
27261 sjöstjärnor 1
27262 sjösäkerhet 4
27263 sjösäkerheten 3
27264 sjösättas 1
27265 sjötransport 1
27266 sjötransporten 1
27267 sjötransporter 3
27268 sjötransportsektorn 1
27269 sjövägen 1
27270 sjövärdighetscertifikat 1
27271 ska 40
27272 skada 38
27273 skadad 1
27274 skadade 6
27275 skadades 2
27276 skadan 3
27277 skadar 17
27278 skadas 2
27279 skadat 3
27280 skadats 6
27281 skadeersättning 1
27282 skadeersättningsanspråk 1
27283 skadeglädje 1
27284 skadegörelse 1
27285 skademinskning 1
27286 skadestånd 1
27287 skadeståndsfrågorna 1
27288 skadlig 8
27289 skadliga 18
27290 skadligare 1
27291 skadligaste 1
27292 skadligt 6
27293 skador 40
27294 skadorna 14
27295 skadornas 2
27296 skaffa 20
27297 skaffade 1
27298 skaffar 2
27299 skaffat 3
27300 skaka 1
27301 skakade 5
27302 skakande 1
27303 skakar 2
27304 skakat 3
27305 skakningar 1
27306 skal 2
27307 skala 7
27308 skalan 1
27309 skaldjur 1
27310 skaldjuren 1
27311 skaldjursfisket 1
27312 skall 1903
27313 skallen 1
27314 skallig 1
27315 skam 7
27316 skamfläck 1
27317 skamlig 3
27318 skamliga 1
27319 skamligt 3
27320 skammen 1
27321 skampålen 3
27322 skandal 7
27323 skandalanklagelserna 1
27324 skandalen 1
27325 skandaler 1
27326 skandalerna 4
27327 skandalös 1
27328 skandalösa 2
27329 skandalöst 5
27330 skapa 292
27331 skapad 1
27332 skapade 9
27333 skapades 6
27334 skapande 7
27335 skapandet 38
27336 skapandets 1
27337 skapar 88
27338 skapare 4
27339 skaparens 1
27340 skaparkraften 1
27341 skapas 44
27342 skapat 22
27343 skapats 20
27344 skapelsen 1
27345 skapelsens 1
27346 skapular 1
27347 skar 2
27348 skara 2
27349 skaran 2
27350 skarp 3
27351 skarpa 4
27352 skarpsinniga 2
27353 skarpt 7
27354 skarv 1
27355 skatt 13
27356 skatta 1
27357 skatte- 2
27358 skatteaspekterna 1
27359 skattebasen 1
27360 skattebestämmelser 1
27361 skattebestämmelserna 1
27362 skattebetalare 10
27363 skattebetalaren 1
27364 skattebetalarna 9
27365 skattebetalarnas 3
27366 skattebördan 1
27367 skatteflykt 1
27368 skattefria 1
27369 skattefrågan 2
27370 skattefrågor 4
27371 skatteförvaltningen 1
27372 skatteförändringar 1
27373 skatteharmonisering 3
27374 skatteharmoniseringen 1
27375 skatteincitament 1
27376 skatteindrivares 1
27377 skatteinkomster 1
27378 skatteinspektörer 1
27379 skattekonkurrens 1
27380 skattelättnader 3
27381 skattemässig 1
27382 skattemässiga 6
27383 skattemässigt 1
27384 skatten 1
27385 skatteområdet 5
27386 skatteparadis 2
27387 skattepengar 2
27388 skattepolitik 3
27389 skattepolitiken 4
27390 skatter 14
27391 skattereform 2
27392 skatteregler 1
27393 skatterna 2
27394 skattesamordning 3
27395 skattesamordningen 1
27396 skattesats 1
27397 skattesatser 1
27398 skattesatserna 1
27399 skattestrukturen 1
27400 skattesystem 2
27401 skattesystemet 4
27402 skattetryck 1
27403 skattetrycket 2
27404 skatteuppgifter 1
27405 skatteändringar 1
27406 skatteåtgärder 1
27407 skattsedeln 2
27408 ske 95
27409 sked 1
27410 skedd 1
27411 skedde 13
27412 skede 17
27413 skeden 1
27414 skedet 2
27415 sken 8
27416 skenat 1
27417 skenet 1
27418 skenhelighet 1
27419 skenheligt 1
27420 skepnader 1
27421 skepp 3
27422 skeppare 1
27423 skeppas 1
27424 skeppat 1
27425 skeppen 1
27426 skeppsbrott 1
27427 skeppsbrottet 1
27428 skeppsbyggnad 1
27429 skeppslanternor 1
27430 skeppsredare 2
27431 skeppsredarnas 1
27432 skeppsvarv 1
27433 skeppsvarven 1
27434 skepsis 2
27435 skepticismen 1
27436 skeptiker 1
27437 skeptisk 6
27438 skeptiska 1
27439 skeptiskt 1
27440 sker 114
27441 skett 49
27442 skick 14
27443 skicka 20
27444 skickad 2
27445 skickade 11
27446 skickades 4
27447 skickar 9
27448 skickas 4
27449 skickat 2
27450 skickats 2
27451 skicklig 3
27452 skicklighet 1
27453 skickligt 2
27454 skifta 2
27455 skiftade 1
27456 skiftande 1
27457 skiftning 1
27458 skikt 2
27459 skilda 14
27460 skilde 1
27461 skildes 2
27462 skildra 1
27463 skildrar 2
27464 skildrats 2
27465 skildring 1
27466 skilja 5
27467 skiljaktigheter 1
27468 skiljaktigheterna 1
27469 skiljas 2
27470 skiljedomare 1
27471 skiljedomarna 1
27472 skiljedomsprövning 1
27473 skiljeförfarandena 1
27474 skiljelinjer 1
27475 skiljer 31
27476 skiljt 1
27477 skillnad 24
27478 skillnaden 13
27479 skillnader 35
27480 skillnaderna 31
27481 skilsmässa 2
27482 skilsmässan 1
27483 skimrade 1
27484 skinande 1
27485 skingra 2
27486 skingrades 1
27487 skinkomeletter 1
27488 skinkor 1
27489 skinkstek 1
27490 skipa 2
27491 skipas 3
27492 skir 1
27493 skiss 3
27494 skissar 1
27495 skissera 3
27496 skisserade 1
27497 skisseras 1
27498 skisserat 2
27499 skit 1
27500 skiva 1
27501 skivor 1
27502 skivsuccéerna 1
27503 skivtallriken 1
27504 skjorta 3
27505 skjortan 3
27506 skjul 3
27507 skjuta 17
27508 skjutas 6
27509 skjutberedd 1
27510 skjuter 9
27511 skjutit 1
27512 skjutits 6
27513 skjuts 9
27514 skjutvapen 1
27515 sko 4
27516 skog 5
27517 skogar 20
27518 skogarna 13
27519 skogarnas 3
27520 skogen 6
27521 skogklädda 1
27522 skogrikedomar 1
27523 skogsarbetarna 1
27524 skogsavverkningen 1
27525 skogsbefolkningens 1
27526 skogsberoende 1
27527 skogsbolagens 1
27528 skogsbruk 1
27529 skogsbrukarna 1
27530 skogsbruket 6
27531 skogsfastighet 1
27532 skogsförordningen 1
27533 skogskommuner 1
27534 skogskornell 1
27535 skogslagar 1
27536 skogsodlingsmaterial 1
27537 skogsområden 1
27538 skogsområdena 1
27539 skogspolitik 1
27540 skogssektorn 3
27541 skogssektorns 1
27542 skogsskövlingen 1
27543 skogsutrustning 1
27544 skogsägaren 2
27545 skojigt 1
27546 skola 7
27547 skolan 9
27548 skolans 1
27549 skolböcker 1
27550 skolelev 1
27551 skolelever 1
27552 skolflickor 1
27553 skollista 1
27554 skolläraraktig 1
27555 skolmaten 1
27556 skolor 4
27557 skolorna 1
27558 skolprefekter 1
27559 skolsalar 1
27560 skolundervisning 1
27561 skolåret 1
27562 skona 2
27563 skonar 1
27564 skonas 1
27565 skoningslös 1
27566 skoningslöst 1
27567 skor 1
27568 skorna 1
27569 skorsten 2
27570 skorstenar 1
27571 skorstenen 1
27572 skotsk 3
27573 skotska 14
27574 skotske 1
27575 skotskt 1
27576 skotten 1
27577 skramlade 1
27578 skrammel 1
27579 skrap 1
27580 skrapa 2
27581 skrapie 11
27582 skrapningar 1
27583 skratt 12
27584 skratta 3
27585 skrattade 12
27586 skrattande 2
27587 skrattas 1
27588 skrattretande 1
27589 skrattspegel 1
27590 skrek 1
27591 skrev 16
27592 skrevs 4
27593 skriade 1
27594 skriande 1
27595 skribenter 1
27596 skrider 1
27597 skriftlig 5
27598 skriftliga 5
27599 skriftligen 8
27600 skriftligt 8
27601 skrik 4
27602 skrika 2
27603 skrikande 1
27604 skrin 1
27605 skriv 1
27606 skriva 24
27607 skrivas 1
27608 skrivberedd 1
27609 skrivbord 1
27610 skrivbordet 1
27611 skrivbordsstolen 1
27612 skrivbordsutvärdering 1
27613 skrivelse 10
27614 skrivelsen 3
27615 skrivelser 2
27616 skriven 2
27617 skriver 9
27618 skrivet 3
27619 skrivit 19
27620 skrivits 2
27621 skrivna 3
27622 skrivningar 1
27623 skrivskyddat 1
27624 skrot 1
27625 skrota 1
27626 skrotade 2
27627 skrotar 2
27628 skrotas 5
27629 skrotfärdigt 1
27630 skrotning 5
27631 skrotningen 2
27632 skrotningsföretag 2
27633 skrotningskostnaden 1
27634 skrotningskostnaderna 1
27635 skrotningsprocesserna 1
27636 skrotningssystem 1
27637 skrov 5
27638 skrovet 2
27639 skrovkonstruktionens 1
27640 skrovsidan 1
27641 skrubb 1
27642 skrubben 2
27643 skrumpnad 1
27644 skrumpnade 1
27645 skrupelfria 2
27646 skrupler 1
27647 skrupulös 1
27648 skrynklade 1
27649 skrynkliga 1
27650 skryt 1
27651 skryta 3
27652 skryter 1
27653 skrytsamt 1
27654 skräck 2
27655 skräckens 1
27656 skräckinjagande 1
27657 skräckscenarior 1
27658 skräckväldet 1
27659 skräddarsydda 1
27660 skräddarsytt 1
27661 skräll 1
27662 skrällande 1
27663 skrämd 1
27664 skrämde 2
27665 skrämma 1
27666 skrämmande 2
27667 skrämmas 1
27668 skrämmer 2
27669 skräms 1
27670 skräp 2
27671 skräpet 2
27672 skräpuppsamlarsyssla 1
27673 skugga 6
27674 skuggad 3
27675 skuggan 4
27676 skuggboxningen 1
27677 skuggig 2
27678 skuggor 2
27679 skuggorna 3
27680 skuggparlament 1
27681 skuld 2
27682 skuldavskrivning 1
27683 skuldbelägger 1
27684 skuldbörda 1
27685 skuldbördan 1
27686 skulden 4
27687 skulder 4
27688 skulderna 1
27689 skuldkvittning 1
27690 skuldmedvetet 1
27691 skuldmedvetna 1
27692 skuldnivåerna 1
27693 skuldnivån 1
27694 skuldsanering 1
27695 skuldsättning 2
27696 skuldsättningen 1
27697 skuldutvecklingen 1
27698 skull 39
27699 skulle 1597
27700 skumma 1
27701 skummjölksblått 1
27702 skumpade 1
27703 skumrasket 1
27704 skumögda 1
27705 skurarna 1
27706 skurits 1
27707 skurkar 1
27708 skurkarna 1
27709 skuta 1
27710 skutan 2
27711 skutt 1
27712 skutta 1
27713 skuttande 1
27714 skvalpade 1
27715 skydd 86
27716 skydda 79
27717 skyddad 1
27718 skyddade 6
27719 skyddande 1
27720 skyddar 12
27721 skyddas 11
27722 skyddat 3
27723 skyddet 49
27724 skydds- 1
27725 skyddsbestämmelser 1
27726 skyddsbestämmelserna 2
27727 skyddsgallren 1
27728 skyddsklausuler 1
27729 skyddslingar 1
27730 skyddslösa 1
27731 skyddsnivå 5
27732 skyddsnivån 4
27733 skyddsnät 2
27734 skyddsnäten 1
27735 skyddsområde 6
27736 skyddsområdet 4
27737 skyddsrum 1
27738 skyddsstyrka 1
27739 skyddssystemen 1
27740 skyddstullar 1
27741 skyddstullarna 1
27742 skyddsvärn 1
27743 skyddsåtgärder 1
27744 skyfall 1
27745 skyfallen 1
27746 skyfflade 1
27747 skygga 1
27748 skygghet 1
27749 skyhöga 1
27750 skyhögt 1
27751 skyla 3
27752 skyldig 14
27753 skyldiga 27
27754 skyldighet 26
27755 skyldigheten 6
27756 skyldigheter 21
27757 skyldigt 2
27758 skylla 1
27759 skyllas 1
27760 skyller 1
27761 skylten 2
27762 skyltfönster 2
27763 skyltfönstret 1
27764 skyltning 1
27765 skymma 2
27766 skymningen 3
27767 skymningsljus 1
27768 skymt 2
27769 skymta 1
27770 skymtade 3
27771 skymtande 2
27772 skymtat 2
27773 skymts 1
27774 skymundan 1
27775 skyn 1
27776 skynda 8
27777 skyndade 3
27778 skyndar 3
27779 skyndsamhet 1
27780 skyndsamt 6
27781 skyttevärn 1
27782 skägget 4
27783 skäggprydd 1
27784 skäggstubb 2
27785 skäl 99
27786 skälen 11
27787 skälet 25
27788 skälig 4
27789 skäliga 4
27790 skäligen 1
27791 skäligt 3
27792 skämdes 1
27793 skämma 1
27794 skämmas 4
27795 skäms 2
27796 skämtar 1
27797 skämtsam 1
27798 skämtsamheter 1
27799 skänka 3
27800 skänker 3
27801 skänkt 2
27802 skänkte 2
27803 skär 7
27804 skära 4
27805 skäras 3
27806 skärmen 5
27807 skärpa 7
27808 skärpas 2
27809 skärper 1
27810 skärpning 2
27811 skärpt 1
27812 skärpta 3
27813 skärrad 1
27814 skärs 2
27815 skärvor 1
27816 skådad 1
27817 skådade 1
27818 skådat 1
27819 skådespel 1
27820 skål 2
27821 skålade 1
27822 skåp 1
27823 skåpdörr 1
27824 skåpet 3
27825 skåra 1
27826 sköldar 1
27827 sköldpaddan 1
27828 skölja 1
27829 sköljde 2
27830 sköna 1
27831 skönhet 6
27832 skönja 1
27833 skönjs 1
27834 skönt 1
27835 skör 1
27836 sköra 2
27837 skörd 3
27838 skörda 1
27839 skördat 1
27840 skörden 1
27841 skörhet 1
27842 sköt 11
27843 sköta 14
27844 skötas 3
27845 sköter 4
27846 sköts 3
27847 skötsamma 1
27848 skötsel 2
27849 skötseln 1
27850 skötselnivå 1
27851 skött 3
27852 skötte 4
27853 skötts 2
27854 skövlade 1
27855 skövling 1
27856 skövlingen 1
27857 slag 45
27858 slagen 1
27859 slaget 7
27860 slagit 10
27861 slagkraftigt 1
27862 slagna 1
27863 slags 60
27864 slak 1
27865 slakt 3
27866 slaktar 2
27867 slaktarna 1
27868 slakten 1
27869 slaktprincip 1
27870 slaktprincipen 1
27871 slam 2
27872 slammer 2
27873 slamrade 1
27874 slamrande 1
27875 slamret 1
27876 slang 1
27877 slank 1
27878 slapp 1
27879 slappa 2
27880 slappare 1
27881 slapphet 5
27882 slappnade 1
27883 slarvigt 1
27884 slav 1
27885 slavar 2
27886 slaveri 2
27887 slem 1
27888 slemmet 1
27889 slemtjockt 1
27890 slet 5
27891 slickade 2
27892 slingor 1
27893 slingrande 3
27894 slint 1
27895 slippa 8
27896 slipper 6
27897 slips 3
27898 slipsen 2
27899 slirar 1
27900 slita 1
27901 sliten 1
27902 sliter 2
27903 slits 1
27904 slitsammaste 1
27905 slockna 2
27906 slocknar 1
27907 slog 28
27908 slogan 1
27909 slogs 2
27910 slokande 1
27911 slopa 2
27912 slopandet 2
27913 slopar 1
27914 slopas 1
27915 slottspark 1
27916 slovenska 1
27917 slovensktalande 1
27918 slug 1
27919 slukade 1
27920 slukar 2
27921 slukas 1
27922 slumområden 1
27923 slump 7
27924 slumpat 1
27925 slumpen 2
27926 slumpmässiga 2
27927 slumpmässigt 1
27928 slumra 1
27929 slumrat 1
27930 slungades 1
27931 slunkit 1
27932 sluppit 1
27933 slussa 1
27934 slussas 1
27935 slut 80
27936 sluta 28
27937 slutade 1
27938 slutande 3
27939 slutandet 1
27940 slutanvändaren 1
27941 slutar 15
27942 slutare 1
27943 slutas 2
27944 slutat 5
27945 slutavtal 1
27946 slutdatum 3
27947 sluten 2
27948 slutenhet 1
27949 sluter 2
27950 slutet 75
27951 slutfasen 1
27952 slutför 1
27953 slutföra 6
27954 slutförande 1
27955 slutförandet 2
27956 slutföras 2
27957 slutförd 1
27958 slutfördes 1
27959 slutförs 2
27960 slutfört 4
27961 slutförts 4
27962 slutgiltig 2
27963 slutgiltiga 15
27964 slutgiltigt 8
27965 sluthanteringen 1
27966 slutit 6
27967 slutits 3
27968 slutkommentar 1
27969 slutkonsumenten 1
27970 slutlig 5
27971 slutliga 23
27972 slutligen 96
27973 slutligt 2
27974 slutmärke 3
27975 slutmärken 1
27976 slutmärkena 1
27977 slutmål 2
27978 slutmålet 1
27979 slutna 4
27980 slutomröstningen 3
27981 slutperioden 1
27982 slutpunkt 2
27983 slutresultat 1
27984 slutresultatet 3
27985 sluts 1
27986 slutsaten 1
27987 slutsats 12
27988 slutsatsen 19
27989 slutsatser 36
27990 slutsatserna 18
27991 slutstatusförhandlingarna 1
27992 sluttning 1
27993 sluttningarna 1
27994 sluttningen 4
27995 slutversionen 1
27996 slutändan 14
27997 slutänden 4
27998 slyngelstater 1
27999 släcka 3
28000 släcker 1
28001 släcks 1
28002 släde 2
28003 släkt 1
28004 släkte 2
28005 släkten 1
28006 släktens 1
28007 släktingar 4
28008 slänga 1
28009 slängde 6
28010 slänger 4
28011 slängs 2
28012 släp 1
28013 släpade 1
28014 släpades 1
28015 släpar 1
28016 släpets 1
28017 släppa 15
28018 släpper 5
28019 släpphänt 1
28020 släpphänta 1
28021 släpphänthet 1
28022 släpphäntheten 2
28023 släppområden 3
28024 släppområdets 1
28025 släppt 1
28026 släppte 6
28027 släpptes 3
28028 släppts 1
28029 släta 2
28030 slätade 1
28031 slätnötta 1
28032 slätt 3
28033 slå 38
28034 slående 1
28035 slår 12
28036 slås 2
28037 slåss 3
28038 slösa 2
28039 slösade 1
28040 slösaktig 1
28041 slösar 1
28042 slösas 4
28043 slösat 1
28044 slösats 1
28045 slöseri 8
28046 slöseriet 1
28047 slöt 4
28048 slöts 1
28049 smak 1
28050 smakar 2
28051 smaken 1
28052 smaklösa 1
28053 smakämnen 1
28054 smal 4
28055 smala 1
28056 smalspårig 1
28057 smalt 1
28058 smekte 1
28059 smickrade 1
28060 smickrar 1
28061 smideskonstens 1
28062 smidig 2
28063 smidigare 1
28064 smidigt 1
28065 smids 1
28066 smita 1
28067 smitning 1
28068 smittad 4
28069 smittade 3
28070 smittades 1
28071 smittar 1
28072 smittas 1
28073 smittsam 2
28074 smittsamma 1
28075 smoking 1
28076 smokingjacka 1
28077 smuggelvaror 1
28078 smugglas 2
28079 smuggling 1
28080 smula 1
28081 smussla 1
28082 smusslande 1
28083 smuts 2
28084 smutsar 1
28085 smutsat 1
28086 smutsbruna 1
28087 smutsig 2
28088 smutsiga 5
28089 smutsigt 2
28090 smycka 1
28091 smycke 1
28092 smyg 1
28093 smyga 2
28094 smygande 1
28095 smyghandlare 1
28096 smäckra 1
28097 smädelse 1
28098 smädelser 1
28099 smäll 2
28100 smälta 3
28101 smältande 1
28102 smärre 2
28103 smärta 6
28104 smärtar 1
28105 smärtas 1
28106 smärtfritt 1
28107 smärtsamma 1
28108 smärtsamt 2
28109 små 125
28110 små- 1
28111 småbarn 2
28112 småbrottslighet 1
28113 småfolket 1
28114 småföretag 8
28115 smågräl 1
28116 småhaiders 1
28117 småhuttra 1
28118 småjordbrukare 1
28119 småningom 14
28120 småpratade 1
28121 småpratar 1
28122 småsak 1
28123 småsaker 2
28124 småskaliga 2
28125 småskaligt 1
28126 småtrevligt 1
28127 smått 1
28128 smög 5
28129 smör 3
28130 smörgås 3
28131 smörgåsar 1
28132 smörgåspaket 1
28133 smörjan 1
28134 smörstekt 1
28135 snabb 19
28136 snabba 24
28137 snabbare 32
28138 snabbast 5
28139 snabbaste 3
28140 snabbhet 2
28141 snabbinsatscentral 1
28142 snabbinsatsstyrka 4
28143 snabbköp 1
28144 snabbt 150
28145 snabbvarningssystem 1
28146 snacka 1
28147 snake-heads 1
28148 snappa 1
28149 snar 10
28150 snarare 62
28151 snarast 30
28152 snaraste 1
28153 snarkade 1
28154 snarlika 1
28155 snart 76
28156 snaskiga 1
28157 snavande 1
28158 sned 1
28159 sneddade 1
28160 snedvrida 2
28161 snedvriden 2
28162 snedvrider 4
28163 snedvridning 12
28164 snedvridningar 6
28165 snedvridningarna 1
28166 snedvridningen 1
28167 snedvridningsriskerna 1
28168 snegla 1
28169 sneglade 1
28170 snett 3
28171 snickra 2
28172 snigeln 3
28173 snigelns 1
28174 snigelpost 1
28175 sniglar 1
28176 snikenhet 1
28177 snikenhetens 1
28178 snirkliga 1
28179 snoriga 1
28180 snubblade 1
28181 snubblande 1
28182 snuddar 1
28183 snurra 2
28184 snurrade 4
28185 snurrar 1
28186 snurrstolar 1
28187 snygg 2
28188 snyggt 1
28189 snäckdjuren 1
28190 snäll 4
28191 snälla 1
28192 snällt 1
28193 snärtar 1
28194 snäste 2
28195 snäv 1
28196 snävare 3
28197 snävt 1
28198 snåren 1
28199 snåriga 1
28200 snöiga 1
28201 snöret 2
28202 snörets 1
28203 snörpvad 2
28204 snörpvadfiske 1
28205 snövit 1
28206 snövitt 1
28207 so 1
28208 social 180
28209 social- 9
28210 sociala 401
28211 socialdemokrater 3
28212 socialdemokraterna 6
28213 socialdemokraternas 3
28214 socialdemokratin 1
28215 socialdemokratisk 3
28216 socialdemokratiska 29
28217 socialdemokratiske 1
28218 socialdemokratiskt 2
28219 socialdepartementet 1
28220 socialekonomisk 1
28221 socialekonomiska 2
28222 socialfonden 14
28223 socialfondens 3
28224 socialfrågor 15
28225 socialförsäkring 1
28226 socialförsäkringen 1
28227 socialförsäkringsfrågor 1
28228 socialförsäkringskostnaderna 1
28229 socialförsäkringsområdet 2
28230 socialförsäkringssystem 3
28231 socialförsäkringssystemen 3
28232 socialhjälp 1
28233 socialist 1
28234 socialister 8
28235 socialisterna 8
28236 socialisternas 1
28237 socialistgruppen 4
28238 socialistgruppens 1
28239 socialistisk 1
28240 socialistiska 19
28241 socialistkollegor 1
28242 socialistparti 1
28243 socialistpartiet 5
28244 socialistpartiets 2
28245 socialministrar 1
28246 socialpolitik 13
28247 socialpolitiken 17
28248 socialpolitikens 1
28249 socialpolitisk 1
28250 socialpolitiska 5
28251 socialrätt 1
28252 socialskyddet 2
28253 socialstatsmodellen 1
28254 socialstöd 3
28255 socialt 61
28256 socialtjänst 1
28257 society 3
28258 socio-ekonomiska 1
28259 socioekonomisk 1
28260 socioekonomiska 6
28261 sociokulturell 1
28262 sociologiska 1
28263 socker 1
28264 sockor 1
28265 sockrat 1
28266 sodomi 1
28267 soffa 1
28268 soffan 4
28269 soffbord 1
28270 soffbordet 1
28271 sofistikerade 2
28272 soft 1
28273 sola 2
28274 solblekta 1
28275 soldaten 1
28276 soldater 15
28277 soldaterna 2
28278 solen 7
28279 solens 1
28280 solglasögon 1
28281 solid 2
28282 solidarisera 1
28283 solidariserade 1
28284 solidarisk 8
28285 solidariska 4
28286 solidariskt 5
28287 solidaritet 62
28288 solidariteten 13
28289 solidaritetens 1
28290 solidaritetsarbetet 1
28291 solidaritetsförhållanden 1
28292 solidaritetssystem 1
28293 solidaritetsuttryck 1
28294 soliditet 1
28295 solig 2
28296 solkant 1
28297 solkungarnas 1
28298 solljus 1
28299 solljuset 3
28300 solnedgången 2
28301 solsken 4
28302 solskenet 3
28303 solstrålarna 1
28304 soluret 1
28305 som 11084
28306 somliga 13
28307 sommar 4
28308 sommaren 12
28309 sommarkvällarna 1
28310 sommarledighet 1
28311 sommarlov 2
28312 sommarlovet 1
28313 sommarnattens 1
28314 sommarsemester 1
28315 somnade 1
28316 son 13
28317 sonen 2
28318 sonens 1
28319 sons 1
28320 sopa 2
28321 sopade 1
28322 sopas 1
28323 sopats 1
28324 soppa 1
28325 sopransångerskor 1
28326 soprantalare 1
28327 soptippen 1
28328 sorg 4
28329 sorgfälligt 1
28330 sorgliga 2
28331 sorgligt 1
28332 sorgsen 1
28333 sorlande 1
28334 sortens 10
28335 sorter 1
28336 sortera 4
28337 sortering 1
28338 sorters 2
28339 sorts 20
28340 sot 4
28341 sotet 1
28342 sov 1
28343 sova 4
28344 sovande 1
28345 sovit 1
28346 sovjetiska 1
28347 sovjettiden 1
28348 sovrummet 4
28349 sovvagn 1
28350 spanjor 6
28351 spanjorer 1
28352 spanjorerna 1
28353 spansk 4
28354 spanska 36
28355 spanske 1
28356 spanskt 2
28357 spara 18
28358 sparade 2
28359 sparande 4
28360 sparandet 1
28361 sparar 4
28362 sparare 1
28363 spararnas 2
28364 sparas 5
28365 sparat 1
28366 sparformer 1
28367 spark 1
28368 sparkar 2
28369 sparkas 1
28370 sparkassor 2
28371 sparmöjligheter 1
28372 sparpengar 2
28373 sparsamma 1
28374 sparvar 1
28375 special 4
28376 specialbestämmelser 4
28377 specialbilaga 1
28378 specialdomstolar 1
28379 specialfiske 1
28380 specialfordon 2
28381 specialförbanden 1
28382 specialinriktning 1
28383 specialiserad 2
28384 specialiserade 4
28385 specialiserat 1
28386 specialiseringen 1
28387 specialister 1
28388 specialistkompetens 1
28389 specialitet 1
28390 specialprogrammen 1
28391 specialtecken 1
28392 specialteckensekvenser 1
28393 specialutbildning 1
28394 speciell 17
28395 speciella 45
28396 speciellt 59
28397 specificera 3
28398 specificerade 1
28399 specificeranden 1
28400 specificerar 2
28401 specificeras 2
28402 specificering 2
28403 specifik 9
28404 specifika 49
28405 specifikation 2
28406 specifikationen 3
28407 specifikationer 1
28408 specifikt 15
28409 speditör 1
28410 speditörerna 1
28411 spegeln 4
28412 spegla 1
28413 speglar 7
28414 speglas 1
28415 speglats 1
28416 spektakel 2
28417 spektakulär 2
28418 spektakulära 1
28419 spektrum 2
28420 spektrumet 3
28421 spekulation 1
28422 spekulationen 1
28423 spekulationer 1
28424 spekulationerna 1
28425 spekulativa 2
28426 spekulativt 1
28427 spekulera 2
28428 spekulerade 1
28429 spel 32
28430 spela 61
28431 spelad 1
28432 spelade 9
28433 spelar 43
28434 spelare 1
28435 spelas 1
28436 spelat 13
28437 spelbrickor 1
28438 spelen 1
28439 spelet 4
28440 spelfält 1
28441 spelfältet 1
28442 spelpjäser 1
28443 spelplan 1
28444 spelregler 8
28445 spelreglerna 2
28446 spelrum 1
28447 spelrummet 1
28448 spendera 3
28449 spenderar 3
28450 spenderas 2
28451 spets 1
28452 spetsade 1
28453 spetsen 6
28454 spetsföretag 1
28455 spetsig 1
28456 spetsiga 2
28457 spettet 1
28458 spika 1
28459 spillo 2
28460 spillolja 2
28461 spillror 1
28462 spills 2
28463 spindelnätet 1
28464 spindlar 1
28465 spionerade 1
28466 spiral 2
28467 spiror 1
28468 spis 1
28469 spisar 1
28470 spisarna 1
28471 spiselhyllan 2
28472 spisen 1
28473 spjut 2
28474 spjutspets 1
28475 split 2
28476 splitterny 1
28477 splittra 1
28478 splittrad 3
28479 splittrade 3
28480 splittras 4
28481 splittrat 2
28482 splittrats 1
28483 splittring 5
28484 spola 1
28485 spolas 2
28486 spongiform 1
28487 sponsorer 1
28488 sponsrad 1
28489 spontan 1
28490 spontana 1
28491 spontaniteten 1
28492 spontant 4
28493 sporadisk 1
28494 sporra 1
28495 sporre 2
28496 sporren 1
28497 sport 1
28498 sportbåtar 1
28499 sportfiskare 1
28500 spots 1
28501 sprack 2
28502 sprang 7
28503 spratt 1
28504 spred 4
28505 spreds 4
28506 spreta 1
28507 spricka 2
28508 sprickan 2
28509 spricker 1
28510 sprickor 1
28511 sprida 9
28512 spridande 1
28513 spridandet 1
28514 spridas 7
28515 spridd 1
28516 spridda 1
28517 sprider 12
28518 spridits 2
28519 spridning 17
28520 spridningen 5
28521 spridningsreglerna 1
28522 sprids 7
28523 springa 5
28524 springande 3
28525 springares 1
28526 springpojke 1
28527 sprit 2
28528 spritts 1
28529 sprudlar 1
28530 sprutade 1
28531 sprutt 1
28532 spräcka 1
28533 sprängande 1
28534 sprängämnen 1
28535 språk 24
28536 språkbruk 3
28537 språken 1
28538 språket 8
28539 språkets 1
28540 språkgrupper 1
28541 språklig 3
28542 språkliga 3
28543 språkområden 1
28544 språkområdena 1
28545 språkversioner 1
28546 språng 2
28547 spurt 1
28548 spy 2
28549 spädbarns 2
28550 spädbarnsdödligheten 1
28551 spänd 3
28552 spända 2
28553 spände 2
28554 spänna 2
28555 spännande 9
28556 spänner 1
28557 spänning 6
28558 spänningar 7
28559 spänningarna 3
28560 spänningen 1
28561 spänningsfält 1
28562 spänningsförhållandet 1
28563 spänst 1
28564 spänt 2
28565 spär 1
28566 spärr 1
28567 spärrar 2
28568 spärras 1
28569 spådomar 1
28570 spår 11
28571 spåra 4
28572 spåras 1
28573 spårbarhet 4
28574 spåren 1
28575 spåret 1
28576 spårning 1
28577 spöke 3
28578 spöken 1
28579 spöklika 1
28580 spökstäder 1
28581 spörsmålet 1
28582 srilankesiska 1
28583 stab 2
28584 stabil 9
28585 stabila 5
28586 stabilare 1
28587 stabilisera 3
28588 stabiliserande 1
28589 stabiliseras 1
28590 stabilisering 4
28591 stabiliseringen 1
28592 stabiliserings- 14
28593 stabiliseringspakten 1
28594 stabiliseringsprocess 1
28595 stabiliseringssträvan 1
28596 stabilitet 38
28597 stabiliteten 15
28598 stabilitetsfaktor 1
28599 stabilitetskursen 1
28600 stabilitetslänk 1
28601 stabilitetspakt 4
28602 stabilitetspakten 20
28603 stabilitetsplanen 1
28604 stabilitetspolitik 1
28605 stabilitetspolitiken 2
28606 stabilt 5
28607 stablitetskultur 1
28608 stack 3
28609 stackars 3
28610 stackatokaskader 1
28611 stad 16
28612 staden 15
28613 stadens 1
28614 stadga 40
28615 stadgan 41
28616 stadgans 1
28617 stadgar 4
28618 stadgehänseende 1
28619 stadier 1
28620 stadiet 3
28621 stadig 2
28622 stadigt 4
28623 stadigvarande 1
28624 stadion 1
28625 stadium 8
28626 stads 1
28627 stads- 2
28628 stadsbefolkningen 1
28629 stadsboende 1
28630 stadsbor 1
28631 stadscentrum 1
28632 stadsdel 1
28633 stadsdelar 2
28634 stadsdelarna 2
28635 stadsdelen 1
28636 stadsförnyelse 1
28637 stadskärnor 2
28638 stadsmiljö 2
28639 stadsmiljögrupp 1
28640 stadsmiljöinitiativ 1
28641 stadsmiljöinitiativet 2
28642 stadsmiljön 1
28643 stadsområde 3
28644 stadsområden 12
28645 stadsområdena 3
28646 stadsområdet 1
28647 stadsplaneringen 1
28648 stadspolitik 1
28649 stadspolitiken 1
28650 stadsrelaterade 1
28651 stadsutveckling 3
28652 stagnation 2
28653 stagnerar 1
28654 stagnerat 2
28655 staka 1
28656 stakeholder 1
28657 stakeholders 1
28658 stalinistiska 1
28659 stalinistiskt 1
28660 stalldörren 1
28661 stammarna 1
28662 stammen 3
28663 stampa 1
28664 stampar 1
28665 stan 5
28666 standard 16
28667 standardanpassningen 1
28668 standarden 2
28669 standarder 8
28670 standardernas 1
28671 standardfilformat 1
28672 standardformatmall 1
28673 standardformuleringar 1
28674 standardfrågeläget 1
28675 standardhöjande 1
28676 standardinställning 1
28677 standardinställningen 1
28678 standardiserade 4
28679 standardiseras 1
28680 standardisering 3
28681 standardiseringar 2
28682 standardiseringen 1
28683 standardiseringskommittén 3
28684 standardiseringssträvandena 2
28685 standards 1
28686 stanna 17
28687 stannade 10
28688 stannande 1
28689 stannar 6
28690 stannat 5
28691 stans 1
28692 staplade 1
28693 stark 43
28694 starka 39
28695 starkare 23
28696 starkast 4
28697 starkaste 5
28698 starke 2
28699 starkt 75
28700 stars 1
28701 start 1
28702 start- 2
28703 start-up-fenomenet 1
28704 start-up-företags 1
28705 starta 16
28706 startade 4
28707 startades 2
28708 startar 4
28709 startas 3
28710 startat 3
28711 startats 3
28712 starten 5
28713 startkapital 1
28714 startmärke 2
28715 startplatta 1
28716 startpunkten 2
28717 stass 1
28718 stat 44
28719 staten 36
28720 statens 9
28721 stater 56
28722 stater-nationer 1
28723 staterna 104
28724 staternas 31
28725 staters 2
28726 station 2
28727 stationen 7
28728 stationens 2
28729 stationerade 1
28730 stationerna 1
28731 stationära 1
28732 statister 1
28733 statistik 14
28734 statistiken 2
28735 statistikens 1
28736 statistisk 3
28737 statistiska 7
28738 statistiskt 4
28739 statlig 11
28740 statliga 75
28741 statligt 28
28742 stats 4
28743 stats- 10
28744 statsbal 1
28745 statsbalen 1
28746 statsbudgeten 1
28747 statschefen 1
28748 statschefer 2
28749 statschefers 1
28750 statsfinanser 1
28751 statsförbund 1
28752 statsgrundandet 1
28753 statskapitalism 1
28754 statskuppen 1
28755 statslösa 1
28756 statsmakt 6
28757 statsmakten 2
28758 statsmaktens 1
28759 statsmakterna 2
28760 statsminister 1
28761 statsministern 1
28762 statsministrarnas 1
28763 statsmonopolet 1
28764 statsmonopolets 1
28765 statsobligationer 1
28766 statssekreteraren 1
28767 statssekreterarens 1
28768 statsskulden 1
28769 statsskulder 1
28770 statsstöd 10
28771 statsstöden 4
28772 statsstödens 3
28773 statsstödet 1
28774 statsstödspolitiken 1
28775 statssäkerheten 1
28776 statstelevision 1
28777 statstjänstemän 1
28778 statsutgifter 1
28779 statsvetare 1
28780 statsvetenskapens 1
28781 statsåklagaren 1
28782 statsöverhuvudena 1
28783 statuera 2
28784 statuerar 1
28785 status 15
28786 statusen 2
28787 stavar 1
28788 stearinljus 2
28789 steering 1
28790 steg 125
28791 stegade 1
28792 stegen 8
28793 steget 8
28794 stegrades 1
28795 stegsumman 1
28796 stegvis 1
28797 stek 1
28798 stekflott 1
28799 stekhus 1
28800 stekpannan 2
28801 stel 3
28802 stela 4
28803 stelt 3
28804 sten 9
28805 stenar 2
28806 stenbeläggning 1
28807 stenbrott 1
28808 stenbyggnader 1
28809 stendövt 1
28810 stenen 1
28811 stenfasaden 1
28812 stenhårda 1
28813 steniga 1
28814 stenigt 1
28815 stenkolen 1
28816 stenkolsindustrierna 1
28817 stenkolsindustrin 2
28818 stenmur 1
28819 stenplattor 1
28820 stereotypa 1
28821 stereotyper 2
28822 steril 1
28823 stetoskopet 1
28824 stick 3
28825 sticka 5
28826 stickande 1
28827 sticker 3
28828 sticket 2
28829 stickord 1
28830 stickprovskontroll 1
28831 stickprovskontroller 1
28832 stickprovstest 1
28833 stickprovsundersökningar 1
28834 stifta 3
28835 stiftar 1
28836 stig 1
28837 stiga 5
28838 stigande 3
28839 stigar 2
28840 stigen 2
28841 stiger 5
28842 stigit 10
28843 stigmatiserat 1
28844 stil 5
28845 stilen 1
28846 stilig 1
28847 stilla 8
28848 stillastående 2
28849 stillhet 3
28850 stillheten 1
28851 stillsamt 2
28852 stimulans 8
28853 stimulansen 3
28854 stimulanser 3
28855 stimulansåtgärder 2
28856 stimulansåtgärderna 1
28857 stimulera 13
28858 stimulerande 7
28859 stimulerar 3
28860 stimulerat 1
28861 stimulering 1
28862 stinkande 1
28863 stint 1
28864 stipulerade 1
28865 stirra 1
28866 stirrade 8
28867 stirrande 1
28868 stirrar 1
28869 stirrat 1
28870 stjäl 1
28871 stjäla 2
28872 stjärna 1
28873 stjärnor 3
28874 stjärnorna 3
28875 stjärnornas 1
28876 stjärt 1
28877 stjärten 1
28878 stockning 1
28879 stocks 1
28880 stod 51
28881 stoft 1
28882 stoftblandning 1
28883 stoftkorn 1
28884 stol 1
28885 stolar 3
28886 stolarna 1
28887 stolen 5
28888 stolsitsen 1
28889 stolt 14
28890 stolta 5
28891 stolte 1
28892 stolthet 8
28893 stoltsera 2
28894 stoltserar 1
28895 stopp 29
28896 stoppa 12
28897 stoppade 3
28898 stoppades 2
28899 stoppar 1
28900 stoppas 9
28901 stoppat 1
28902 stoppats 1
28903 stor 306
28904 stora 347
28905 storartad 1
28906 storartat 2
28907 stordrifts- 1
28908 stordriftsfördelar 1
28909 stordriftsfördelarna 1
28910 store 1
28911 storföretag 2
28912 storföretagens 1
28913 storhet 2
28914 storheter 1
28915 storhetsvansinne 1
28916 storkapitalet 1
28917 storkapitalets 2
28918 storkonsument 1
28919 storlek 6
28920 storleken 4
28921 storleksordningen 3
28922 storm 2
28923 stormakt 1
28924 stormakterna 1
28925 stormar 7
28926 stormarknader 2
28927 stormarna 12
28928 stormarnas 1
28929 stormen 6
28930 stormens 1
28931 stormfloden 1
28932 stormfällda 1
28933 stormvind 1
28934 storsinta 1
28935 storskalig 1
28936 storskaliga 4
28937 storskalighet 1
28938 storslaget 1
28939 storslagna 2
28940 storstadsförorter 1
28941 storstäderna 3
28942 stort 132
28943 stortårna 1
28944 storvulen 1
28945 straff 10
28946 straff- 2
28947 straffa 4
28948 straffas 3
28949 straffats 1
28950 straffbar 2
28951 straffbara 1
28952 straffbarheten 1
28953 straffbart 1
28954 straffbestämmelser 1
28955 straffet 2
28956 strafflagstiftning 2
28957 straffläger 1
28958 strafflöshet 1
28959 straffprocessrätten 1
28960 straffprocessrättsligt 1
28961 straffrihet 1
28962 straffriheten 1
28963 straffrätt 10
28964 straffrätten 12
28965 straffrättens 3
28966 straffrättslig 3
28967 straffrättsliga 32
28968 straffrättsligt 10
28969 straffrättsområdet 1
28970 stram 3
28971 strama 2
28972 stramhet 1
28973 strand 1
28974 stranda 1
28975 stranden 4
28976 strandremsa 4
28977 strandremsan 2
28978 strandremsans 1
28979 strategi 86
28980 strategidokument 2
28981 strategier 37
28982 strategierna 3
28983 strategin 19
28984 strategiplanering 1
28985 strategisk 11
28986 strategiska 51
28987 strategiskt 13
28988 strax 13
28989 strecksats 1
28990 stress 1
28991 stretar 1
28992 strid 24
28993 strida 6
28994 stridande 1
28995 striden 3
28996 strider 25
28997 stridigheten 1
28998 stridsropet 1
28999 stridsvagnar 1
29000 strikt 25
29001 strikta 17
29002 striktare 6
29003 strimma 2
29004 strimman 1
29005 strimmorna 1
29006 stringens 1
29007 stringentare 1
29008 stripes 1
29009 stripigt 1
29010 strukits 2
29011 struktur 32
29012 strukturanpassningen 1
29013 strukturell 7
29014 strukturella 25
29015 strukturellt 6
29016 strukturen 17
29017 strukturer 34
29018 strukturera 1
29019 strukturerad 3
29020 strukturerande 2
29021 strukturerar 1
29022 struktureras 1
29023 strukturerat 6
29024 struktureringen 1
29025 strukturerna 8
29026 strukturers 1
29027 strukturfonden 3
29028 strukturfonder 18
29029 strukturfonderna 96
29030 strukturfonderna- 1
29031 strukturfondernas 6
29032 strukturfondsmedel 1
29033 strukturfondsprogram 1
29034 strukturfondsprogrammen 2
29035 strukturfondsrunda 1
29036 strukturfondsstödet 1
29037 strukturformerna 2
29038 strukturförändringen 1
29039 strukturmässig 1
29040 strukturpolitik 8
29041 strukturpolitiken 5
29042 strukturprojekt 1
29043 strukturreformer 3
29044 strukturstramhet 1
29045 strukturstöd 4
29046 strukturstöden 1
29047 strukturutgifterna 1
29048 strukturutveckling 2
29049 strukturåtgärderna 1
29050 strumpor 2
29051 strumporna 1
29052 strumpstickor 1
29053 strumpsömmar 1
29054 strunta 5
29055 struntar 3
29056 struntat 1
29057 struntprat 3
29058 strupen 1
29059 struts 1
29060 stryk 1
29061 stryka 5
29062 strykas 2
29063 strykningen 1
29064 stryks 3
29065 stryps 1
29066 strypt 1
29067 sträck 1
29068 sträcka 9
29069 sträckan 1
29070 sträcker 9
29071 sträckor 1
29072 sträckte 5
29073 stränder 10
29074 stränderna 6
29075 sträng 8
29076 stränga 14
29077 strängare 5
29078 strängaste 2
29079 stränghet 4
29080 strängt 9
29081 sträva 16
29082 strävade 2
29083 strävan 27
29084 strävanden 7
29085 strävandena 1
29086 strävar 20
29087 strävat 1
29088 strået 2
29089 strålande 2
29090 strålar 1
29091 stråle 1
29092 strålkastare 1
29093 strålkastaren 1
29094 strålkastarljuset 1
29095 strålning 1
29096 strålskydd 1
29097 strödde 1
29098 strök 1
29099 ströks 1
29100 ström 5
29101 strömmade 3
29102 strömmande 2
29103 strömmarna 1
29104 strömningar 4
29105 strömningarna 1
29106 strömningen 2
29107 ströva 1
29108 strövade 1
29109 stuckit 1
29110 student 3
29111 studenten 1
29112 studenter 3
29113 studenterna 1
29114 studentskan 1
29115 studera 2
29116 studerade 2
29117 studerar 4
29118 studeras 2
29119 studerat 3
29120 studie 6
29121 studiebesök 1
29122 studiedag 1
29123 studien 1
29124 studieprogram 1
29125 studier 16
29126 studsade 2
29127 stugor 1
29128 stum 3
29129 stund 31
29130 stundande 3
29131 stunden 3
29132 stunder 4
29133 stunderna 1
29134 stundtals 1
29135 stuvade 1
29136 stycke 4
29137 stycken 3
29138 styckena 2
29139 stycket 4
29140 stympad 2
29141 stympningen 1
29142 styr 6
29143 styra 19
29144 styrande 2
29145 styras 6
29146 styrd 1
29147 styrda 1
29148 styrde 4
29149 styre 3
29150 styrekonomen 3
29151 styrelse 3
29152 styrelsebeslut 1
29153 styrelseformer 1
29154 styrelseformerna 1
29155 styrelsen 3
29156 styrelser 1
29157 styrelseskick 1
29158 styret 2
29159 styrets 1
29160 styrka 13
29161 styrkan 4
29162 styrkeförhållandena 2
29163 styrkeposition 1
29164 styrketest 1
29165 styrkommittéerna 1
29166 styrkor 15
29167 styrkorna 5
29168 styrning 2
29169 styrningen 2
29170 styrs 5
29171 styrt 3
29172 styva 1
29173 styvsint 1
29174 styvt 1
29175 städ 1
29176 städa 5
29177 städade 2
29178 städat 1
29179 städer 27
29180 städerna 27
29181 städernas 5
29182 städers 2
29183 städning 1
29184 ställ 1
29185 ställa 95
29186 ställas 32
29187 ställda 2
29188 ställde 28
29189 ställdes 6
29190 ställe 15
29191 ställen 9
29192 ställer 68
29193 stället 135
29194 ställning 73
29195 ställningar 1
29196 ställningen 1
29197 ställningstagande 12
29198 ställningstaganden 4
29199 ställningstagandet 1
29200 ställs 30
29201 ställt 24
29202 ställts 8
29203 stämde 3
29204 stämma 6
29205 stämmer 35
29206 stämning 1
29207 stämningen 3
29208 stämningsansökningar 1
29209 stämpling 1
29210 ständig 7
29211 ständiga 15
29212 ständigt 45
29213 stänga 3
29214 stängda 2
29215 stängde 4
29216 stänger 3
29217 stängerna 1
29218 stängning 3
29219 stängningen 2
29220 stängs 3
29221 stängsel 1
29222 stängts 3
29223 stänkte 1
29224 stärka 65
29225 stärkande 6
29226 stärkandet 4
29227 stärkas 8
29228 stärker 9
29229 stärks 5
29230 stärkt 3
29231 stärkts 2
29232 stäv 3
29233 stävja 1
29234 stävjas 1
29235 stå 66
29236 stående 7
29237 stål 1
29238 stålföretag 5
29239 stålgemenskapen 1
29240 stålindustrin 23
29241 stålindustrins 2
29242 stålsektorn 4
29243 stålverk 2
29244 stålverket 2
29245 stålverksanläggningar 1
29246 stånd 60
29247 ståndpunkt 137
29248 ståndpunkten 65
29249 ståndpunkter 41
29250 ståndpunkterna 5
29251 ståndpunktstagande 1
29252 stång 1
29253 står 254
29254 ståtlig 2
29255 stått 18
29256 stöd 344
29257 stöd- 1
29258 stödbehov 1
29259 stödberättigade 7
29260 stödberättigande 1
29261 stödd 3
29262 stödda 1
29263 stödde 6
29264 stöddes 1
29265 stöden 26
29266 stöder 162
29267 stödet 51
29268 stödets 1
29269 stödformer 1
29270 stödinstrument 1
29271 stödja 165
29272 stödjande 3
29273 stödjas 14
29274 stödjer 5
29275 stödkategorier 1
29276 stödköper 1
29277 stödmedlen 1
29278 stödmekanismer 1
29279 stödmottagaren 1
29280 stödmöjligheter 1
29281 stödnivån 2
29282 stödområden 1
29283 stödområdena 1
29284 stödpolitik 1
29285 stödprogram 5
29286 stödpunkt 1
29287 stödpunkten 1
29288 stödram 1
29289 stödramar 1
29290 stöds 16
29291 stödsystem 3
29292 stödsystemet 1
29293 stödsänkningarna 1
29294 stödverktygen 1
29295 stödyta 1
29296 stödåtgärder 11
29297 stödåtgärderna 2
29298 stöld 3
29299 stönade 1
29300 stöpa 2
29301 stöpsleven 1
29302 stör 4
29303 störa 3
29304 störande 3
29305 störas 1
29306 störd 1
29307 störde 2
29308 störning 1
29309 störningar 5
29310 störningarna 1
29311 större 207
29312 störs 2
29313 störst 9
29314 största 103
29315 störste 1
29316 störta 3
29317 störtade 2
29318 störtflod 1
29319 stöt 3
29320 stöta 2
29321 stötande 1
29322 stöten 1
29323 stöter 2
29324 stötestenarna 1
29325 stötfångare 1
29326 stött 19
29327 stötta 2
29328 stöttat 2
29329 stötte 5
29330 stöttepelare 1
29331 stöttepelaren 1
29332 stötts 2
29333 sua 1
29334 sub 1
29335 subject 1
29336 subjekt 1
29337 subjektiva 1
29338 sublima 1
29339 subsidaritetsprincipen 2
29340 subsidiaritet 10
29341 subsidiariteten 11
29342 subsidiaritets- 1
29343 subsidiaritetsaltaret 1
29344 subsidiaritetsfrågor 2
29345 subsidiaritetsprincip 1
29346 subsidiaritetsprincipen 28
29347 subsidiaritetsprinciper 1
29348 subsidiär 1
29349 substans 2
29350 substansen 1
29351 substantiella 2
29352 substantiellt 1
29353 substitut 2
29354 subtila 1
29355 subvention 1
29356 subventioner 12
29357 subventionera 3
29358 subventionerade 1
29359 subventionerar 1
29360 subventioneras 1
29361 subventionerna 2
29362 subventionskonkurrens 1
29363 successiv 2
29364 successiva 4
29365 successivt 7
29366 suckade 1
29367 suckades 1
29368 sudaneserna 1
29369 sudda 2
29370 suddades 1
29371 suddig 1
29372 suger 1
29373 sugs 1
29374 summa 6
29375 summan 2
29376 summarisk 1
29377 summera 1
29378 summertonen 1
29379 summor 13
29380 sund 4
29381 sunda 7
29382 sundare 3
29383 sundaste 1
29384 sundhet 1
29385 sunt 4
29386 supa 1
29387 supereuropéerna 1
29388 supermakt 2
29389 superstat 1
29390 supranationell 1
29391 surrad 1
29392 surrogat 1
29393 surrogatfader 2
29394 surögt 1
29395 susade 1
29396 suspekta 1
29397 suspenderas 1
29398 suspensiv 1
29399 suttit 7
29400 suverän 2
29401 suveräna 5
29402 suveränitet 19
29403 suveräniteten 6
29404 suveränt 1
29405 svag 11
29406 svaga 12
29407 svagare 10
29408 svagares 1
29409 svagaste 5
29410 svaghet 11
29411 svagheten 3
29412 svagheter 4
29413 svagheterna 3
29414 svagt 3
29415 svaj 1
29416 svajade 1
29417 sval 1
29418 svalde 1
29419 svansar 1
29420 svansen 1
29421 svar 121
29422 svara 44
29423 svarade 22
29424 svarande 1
29425 svarar 17
29426 svarat 8
29427 svaren 7
29428 svaret 25
29429 svaromål 1
29430 svars 9
29431 svarstider 1
29432 svarston 1
29433 svart 17
29434 svarta 15
29435 svartas 1
29436 svarte 1
29437 svartingar 2
29438 svartingarna 1
29439 svartjobb 1
29440 svartklädda 2
29441 svartkonst 1
29442 svartkonstnären 1
29443 svartlista 1
29444 svartröd 1
29445 svassa 1
29446 svavelhalt 1
29447 svavelhalten 1
29448 svek 3
29449 svekfullt 1
29450 svensk 4
29451 svenska 22
29452 svenskarna 1
29453 svenske 1
29454 svensken 1
29455 svenskt 1
29456 svepande 1
29457 svepskäl 2
29458 svepte 3
29459 svett 2
29460 svetten 2
29461 svettglänsande 1
29462 svikit 1
29463 svinaktigt 1
29464 svindel 2
29465 svindlande 1
29466 svinstia 1
29467 svischade 1
29468 sviterna 1
29469 svurit 1
29470 svällande 1
29471 svält 4
29472 svältsituationer 1
29473 svämmade 1
29474 svämmar 1
29475 svänga 1
29476 svängande 1
29477 svängd 1
29478 svängde 4
29479 svängningar 1
29480 svängrum 1
29481 svär 1
29482 svärd 1
29483 svärdet 1
29484 svärta 2
29485 svärtas 1
29486 sväva 1
29487 svävade 3
29488 svävande 4
29489 svåger 1
29490 svågerpolitik 3
29491 svål 1
29492 svångrems- 1
29493 svår 28
29494 svåra 45
29495 svårare 10
29496 svårartade 1
29497 svåraste 2
29498 svårbedömbara 1
29499 svårbegriplig 2
29500 svårhanterliga 1
29501 svårighet 2
29502 svårigheten 3
29503 svårigheter 69
29504 svårigheterna 13
29505 svårligen 1
29506 svårlöst 1
29507 svårlösta 1
29508 svårmod 1
29509 svårt 96
29510 svårtolkat 1
29511 svåröverskådligt 1
29512 svåröverstigliga 1
29513 syd 1
29514 sydafrikanen 2
29515 sydafrikanens 1
29516 sydafrikanerna 1
29517 sydafrikanska 1
29518 sydamerikanska 1
29519 sydeuropeiska 1
29520 sydkusten 1
29521 sydlig 1
29522 sydliga 2
29523 sydligt 1
29524 sydvästra 2
29525 sydöstra 10
29526 syfta 2
29527 syftade 5
29528 syftande 1
29529 syftar 79
29530 syfte 85
29531 syften 13
29532 syftena 2
29533 syftet 40
29534 sykomorträ 1
29535 symbol 8
29536 symbolen 1
29537 symboler 1
29538 symbolerna 1
29539 symbolisera 1
29540 symboliserar 1
29541 symbolisk 5
29542 symboliska 4
29543 symboliskt 1
29544 symbolism 1
29545 symfoniorkestrar 1
29546 sympati 10
29547 sympatier 1
29548 sympatiserade 1
29549 sympatiserar 3
29550 sympatiskt 2
29551 sympatiyttring 1
29552 symptom 3
29553 symptomatiska 1
29554 symptomen 1
29555 symtom 2
29556 syn 31
29557 syna 1
29558 synar 1
29559 synas 3
29560 synd 11
29561 syndabock 1
29562 syndabockar 2
29563 syndar 1
29564 synder 1
29565 syndikalister 2
29566 syndromet 1
29567 synen 3
29568 synergi 1
29569 synergieffekter 3
29570 synergierna 1
29571 synergism 1
29572 synes 4
29573 synfält 1
29574 synhåll 2
29575 synkroniserad 1
29576 synkroniseringen 1
29577 synlig 5
29578 synliga 6
29579 synligare 1
29580 synligaste 1
29581 synliggörs 1
29582 synligt 2
29583 synnerhet 163
29584 synnerligen 17
29585 synonym 1
29586 synonymt 1
29587 synpunkt 18
29588 synpunkten 7
29589 synpunkter 47
29590 synpunkterna 2
29591 syns 2
29592 synsätt 13
29593 synsättet 1
29594 syntax-regler 1
29595 syntes 5
29596 syntetiska 1
29597 synvinkel 26
29598 synvinkeln 8
29599 synvinklar 1
29600 syrier 1
29601 syrierna 3
29602 syriska 4
29603 syriske 1
29604 sysselsatt 3
29605 sysselsatta 3
29606 sysselsätta 2
29607 sysselsätter 4
29608 sysselsättning 195
29609 sysselsättningen 87
29610 sysselsättningens 3
29611 sysselsättnings- 3
29612 sysselsättningsargumentet 1
29613 sysselsättningsbas 1
29614 sysselsättningsdrivande 1
29615 sysselsättningsfaktor 1
29616 sysselsättningsfluktuationerna 1
29617 sysselsättningsfrämjande 2
29618 sysselsättningsfrågan 2
29619 sysselsättningsförhållanden 1
29620 sysselsättningsförmåga 3
29621 sysselsättningsgrad 4
29622 sysselsättningsinitiativ 1
29623 sysselsättningsinitiativen 1
29624 sysselsättningskvaliteten 1
29625 sysselsättningsläget 1
29626 sysselsättningsmodeller 1
29627 sysselsättningsmöjligheter 2
29628 sysselsättningsnivå 4
29629 sysselsättningsnivåer 1
29630 sysselsättningsnivåerna 1
29631 sysselsättningsnivån 4
29632 sysselsättningsområden 1
29633 sysselsättningsområdet 2
29634 sysselsättningspaketet 1
29635 sysselsättningspakten 1
29636 sysselsättningspakterna 1
29637 sysselsättningsplaner 1
29638 sysselsättningspolitik 11
29639 sysselsättningspolitiken 15
29640 sysselsättningspolitiska 6
29641 sysselsättningspotential 2
29642 sysselsättningsproblem 2
29643 sysselsättningsproblematiken 2
29644 sysselsättningsprogrammen 1
29645 sysselsättningsrapporten 2
29646 sysselsättningssamarbetet 1
29647 sysselsättningsskapande 6
29648 sysselsättningsskydd 1
29649 sysselsättningsstrategi 2
29650 sysselsättningsstrategier 1
29651 sysselsättningsstrategin 7
29652 sysselsättningsstrategins 1
29653 sysselsättningstoppmötet 1
29654 sysselsättningsvänliga 1
29655 sysselsättningsåtgärder 1
29656 sysselsättningsåtgärderna 1
29657 sysselsättningsökningen 1
29658 syssla 3
29659 sysslade 3
29660 sysslar 9
29661 sysslolösa 3
29662 system 173
29663 systematisera 1
29664 systematisk 10
29665 systematiska 2
29666 systematiskt 12
29667 systemen 20
29668 systemet 78
29669 systemets 1
29670 systemmodernisering 1
29671 systemutveckling 1
29672 systemändring 2
29673 systemändringen 1
29674 syster 3
29675 systerfartyg 1
29676 systern 1
29677 systerskap 1
29678 systerson 1
29679 systrar 4
29680 säden 1
29681 säg 2
29682 säga 529
29683 sägas 12
29684 säger 235
29685 sägs 17
29686 säker 69
29687 säkerhet 140
29688 säkerheten 48
29689 säkerhetens 2
29690 säkerhets 2
29691 säkerhets- 8
29692 säkerhetsanordning 1
29693 säkerhetsargument 1
29694 säkerhetsaspekten 1
29695 säkerhetsbestämmelser 2
29696 säkerhetsbestämmelserna 1
29697 säkerhetsbältet 1
29698 säkerhetsfrågan 2
29699 säkerhetsfrågor 2
29700 säkerhetsfångar 1
29701 säkerhetsföreskrifterna 1
29702 säkerhetsförhållandena 1
29703 säkerhetsgarantierna 2
29704 säkerhetsgränsen 1
29705 säkerhetshänsyn 1
29706 säkerhetsinsatserna 1
29707 säkerhetsinställningar 1
29708 säkerhetsintresse 1
29709 säkerhetskontrollerna 1
29710 säkerhetskopia 1
29711 säkerhetskopian 1
29712 säkerhetskriser 1
29713 säkerhetsnivå 1
29714 säkerhetsnivån 1
29715 säkerhetsnormer 2
29716 säkerhetsnätet 1
29717 säkerhetsorganisation 1
29718 säkerhetspolitik 15
29719 säkerhetspolitiken 8
29720 säkerhetspolitikens 1
29721 säkerhetspolitisk 1
29722 säkerhetsproblem 2
29723 säkerhetsproblemen 1
29724 säkerhetsrisk 3
29725 säkerhetsrisker 1
29726 säkerhetsråd 7
29727 säkerhetsrådet 2
29728 säkerhetsrådets 4
29729 säkerhetsrådgivare 12
29730 säkerhetsrådgivarna 1
29731 säkerhetsråds 1
29732 säkerhetsskäl 1
29733 säkerhetsstyrka 1
29734 säkerhetsstyrkans 1
29735 säkerhetsställande 1
29736 säkerhetssystemet 1
29737 säkerhetstjänst 1
29738 säkerhetsventil 1
29739 säkerhetsåtgärd 1
29740 säkerhetsåtgärderna 1
29741 säkerhetsövningar 1
29742 säkerligen 22
29743 säkerställa 55
29744 säkerställande 1
29745 säkerställandet 2
29746 säkerställas 1
29747 säkerställd 1
29748 säkerställer 12
29749 säkerställs 1
29750 säkerställt 1
29751 säkert 60
29752 säkerthetsnormer 1
29753 säkra 43
29754 säkrad 3
29755 säkrade 2
29756 säkrandet 3
29757 säkrar 3
29758 säkrare 4
29759 säkras 3
29760 säkraste 5
29761 säkrat 1
29762 sälja 10
29763 säljare 3
29764 säljas 7
29765 säljer 4
29766 säljförbud 1
29767 säljs 1
29768 säljstart 1
29769 sällan 9
29770 sällsamheter 1
29771 sällsamma 1
29772 sällskap 5
29773 sällskapliga 1
29774 sällskaplighet 1
29775 sällsynt 3
29776 sämre 20
29777 sämst 8
29778 sämsta 1
29779 sända 12
29780 sändas 3
29781 sände 3
29782 sändebud 9
29783 sändebudet 4
29784 sänder 3
29785 sändes 1
29786 sändningar 1
29787 sändningarna 1
29788 sändningsläge 1
29789 sänds 3
29790 säng 2
29791 sängen 5
29792 sängkammare 1
29793 sängkläderna 1
29794 sängs 1
29795 sänka 14
29796 sänkan 1
29797 sänkas 3
29798 sänker 1
29799 sänkning 3
29800 sänkningar 1
29801 sänkningen 2
29802 sänks 1
29803 sänkt 1
29804 sänkta 1
29805 sänkte 2
29806 sänkts 1
29807 sänt 2
29808 sär 1
29809 särart 1
29810 särarten 1
29811 särarter 1
29812 särbehandla 1
29813 särbehandling 6
29814 särbestämmelse 1
29815 särbestämmelser 1
29816 särdrag 9
29817 särdragen 1
29818 säreget 1
29819 säregna 1
29820 särintressen 2
29821 särkilt 1
29822 särskild 44
29823 särskilda 54
29824 särskilja 2
29825 särskilt 377
29826 säsong 2
29827 säsongsarbete 1
29828 säsongsarbetslöshet 1
29829 säsongsbetonad 1
29830 säsongsbetonade 1
29831 säsongsbundna 2
29832 säsongsjobb 1
29833 säte 4
29834 säten 1
29835 sätet 2
29836 sätt 684
29837 sätta 91
29838 sättandes 1
29839 sättas 14
29840 sätten 3
29841 sätter 34
29842 sättet 71
29843 sätts 14
29844 sättstycken 1
29845 sävliga 1
29846 så 1741
29847 sådan 196
29848 sådana 139
29849 sådant 145
29850 såg 89
29851 såga 1
29852 sågs 1
29853 sågspån 1
29854 sågverk 1
29855 såhär 2
29856 sålde 4
29857 såldes 1
29858 således 131
29859 såll 3
29860 sållas 1
29861 sålt 1
29862 sålts 1
29863 sålunda 10
29864 sån 8
29865 såna 5
29866 sång 1
29867 sången 1
29868 sångens 1
29869 sånger 1
29870 sånt 2
29871 såra 1
29872 sårade 2
29873 sårbar 1
29874 sårbara 8
29875 sårbarhet 1
29876 sårbarheten 1
29877 såsom 103
29878 såtillvida 2
29879 såvida 7
29880 såvitt 2
29881 såväl 122
29882 söder 23
29883 söderut 2
29884 södra 26
29885 sögs 1
29886 söka 15
29887 sökande 4
29888 sökanden 1
29889 sökandet 4
29890 sökas 2
29891 söker 24
29892 sökningen 1
29893 sökt 1
29894 sökte 5
29895 sökväg 5
29896 sökvägen 1
29897 sömn 2
29898 söndags 1
29899 söndagstidningar 1
29900 sönder 9
29901 sönderdela 2
29902 sönderdelas 1
29903 sönderdelning 1
29904 sönderdelningsanläggningarna 1
29905 sönderfall 2
29906 söndergrävd 1
29907 sönderklippta 1
29908 sönderrivna 1
29909 sönderslaget 1
29910 sönderslagna 1
29911 söner 4
29912 sörja 10
29913 sörjde 2
29914 sörjer 6
29915 söt 1
29916 sötvatten 1
29917 sötvattenmatros 1
29918 t 2
29919 t. 1
29920 t.ex 6
29921 t.ex. 59
29922 t.o.m. 18
29923 ta 643
29924 tabell 5
29925 tabellen 3
29926 tabeller 5
29927 tabellerna 2
29928 tabletter 1
29929 tabu 1
29930 tabubelagda 1
29931 tabubelagt 1
29932 tack 91
29933 tacka 178
29934 tackar 58
29935 tacklas 1
29936 tacknämligt 2
29937 tackor 1
29938 tacksam 23
29939 tacksamhet 2
29940 tacksamhetens 1
29941 tacksamma 5
29942 tacksamt 1
29943 tag 14
29944 tagen 3
29945 taget 55
29946 tagit 117
29947 tagits 36
29948 tagna 2
29949 tak 8
29950 taken 1
29951 taket 11
29952 takt 14
29953 takten 5
29954 takter 1
29955 taktik 7
29956 taktiska 2
29957 taktiskt 1
29958 taktlöshet 1
29959 takåsarna 1
29960 tal 50
29961 tala 158
29962 talade 79
29963 talades 3
29964 talan 3
29965 talande 1
29966 talang 1
29967 talanger 2
29968 talar 157
29969 talare 36
29970 talaren 11
29971 talares 1
29972 talarlistan 1
29973 talarna 13
29974 talarnas 1
29975 talarstolen 1
29976 talartid 5
29977 talartiden 3
29978 talartiderna 2
29979 talas 28
29980 talat 48
29981 talats 2
29982 talen 2
29983 talesman 5
29984 talesmannen 1
29985 talesmän 1
29986 talesätt 1
29987 talesättet 1
29988 talet 6
29989 talförmågan 1
29990 tallitkatan 1
29991 tallrik 4
29992 tallrikar 1
29993 tallrikarna 1
29994 tallriken 3
29995 tallöst 1
29996 talman 1137
29997 talmannen 11
29998 talmannens 2
29999 talmans 2
30000 talmanskonferens 1
30001 talmanskonferensen 15
30002 talmanskonferenser 1
30003 talmän 2
30004 talrika 6
30005 tals 3
30006 tampas 2
30007 tandem 1
30008 tandlöst 1
30009 tangera 1
30010 tank- 1
30011 tankar 32
30012 tankarna 14
30013 tankbåtar 1
30014 tankbåtarna 2
30015 tanke 151
30016 tankearbetet 1
30017 tankebanor 1
30018 tankefrihet 1
30019 tankegångar 2
30020 tankegångarna 2
30021 tankemöda 1
30022 tanken 40
30023 tankens 1
30024 tankepolis 1
30025 tankern 1
30026 tankerägarnas 1
30027 tankespår 1
30028 tankfartyg 7
30029 tankfartygens 1
30030 tankfartyget 3
30031 tankfordon 1
30032 tankfull 1
30033 tanklöshet 1
30034 tanklöst 1
30035 tankrengöring 2
30036 tankrengöringar 1
30037 tankrengöringarna 1
30038 tapeten 1
30039 tappa 6
30040 tappar 3
30041 tappat 2
30042 tappert 1
30043 tappt 1
30044 tar 219
30045 tarifferna 1
30046 tarvligheter 2
30047 tas 131
30048 task 1
30049 tatuerat 1
30050 tavlor 2
30051 tavlorna 1
30052 tax-free 1
30053 tax-free-försäljningen 1
30054 tax-free-lobbyister 1
30055 taxa 1
30056 taxeringsnormer 1
30057 taxi 3
30058 taxichaufför 1
30059 taxifolia 1
30060 taxin 2
30061 taxor 1
30062 taxorna 1
30063 tayloristiska 1
30064 te 1
30065 teater 1
30066 teaterföreställning 1
30067 teatergrupper 1
30068 tecken 26
30069 tecknade 1
30070 tecknas 1
30071 tecknats 1
30072 tecknen 1
30073 tedde 2
30074 tegel 2
30075 tegeldamm 1
30076 tegelskärva 1
30077 teknik 24
30078 tekniken 16
30079 teknikens 2
30080 tekniker 8
30081 teknikerna 6
30082 teknisk 38
30083 teknisk-ekonomiskt 1
30084 tekniska 86
30085 tekniskt 26
30086 teknokraternas 1
30087 teknologi 3
30088 teknologiska 1
30089 telefon 5
30090 telefonavlyssning 4
30091 telefonavlyssningen 1
30092 telefonbolaget 1
30093 telefonen 2
30094 telefoner 1
30095 telefoni 1
30096 telefonicentren 1
30097 telefonisterna 1
30098 telefonitjänster 1
30099 telefonnummer 1
30100 telefonsamtal 3
30101 telefonsamtalet 1
30102 teleföretagen 1
30103 telegram 2
30104 telekommunikation 4
30105 telekommunikationen 1
30106 telekommunikationer 2
30107 telekommunikationernas 1
30108 telekommunikationsministern 1
30109 telekommunikationsområdet 1
30110 telekommunikationspriserna 1
30111 telekommunikationssektorn 1
30112 telenät 1
30113 teletrafiken 2
30114 televerket 1
30115 television 1
30116 televisionen 3
30117 televisionsprogrammen 1
30118 tema 1
30119 temat 1
30120 tematisk 2
30121 tematiska 4
30122 tempel 1
30123 temperatur 2
30124 temperaturen 3
30125 temperaturer 4
30126 temperaturhöjningar 1
30127 tempererad 1
30128 tempo 3
30129 temporär 2
30130 temporärt 1
30131 tempot 1
30132 tendens 11
30133 tendensen 9
30134 tendenser 2
30135 tendenserna 3
30136 tendentiöst 1
30137 tenderar 9
30138 tennisbollar 1
30139 teokratiskt 1
30140 teologerna 1
30141 teologi 1
30142 teoretisk 2
30143 teoretiska 2
30144 teoretiskt 7
30145 teori 3
30146 teorier 1
30147 teorin 4
30148 ter 1
30149 teratogena 1
30150 teratogent 1
30151 term 2
30152 termen 3
30153 termer 9
30154 termerna 1
30155 terminaler 1
30156 terminen 1
30157 terminis 2
30158 terminologi 1
30159 termins- 1
30160 terminskontrakt 2
30161 territorialitetsprincipen 1
30162 territorialklausul 1
30163 territorialklausulen 3
30164 territorialvatten 1
30165 territorieklausulen 1
30166 territoriell 2
30167 territoriella 15
30168 territorier 5
30169 territoriet 7
30170 territoriets 1
30171 territorium 30
30172 terror 1
30173 terrorbomb 1
30174 terrorism 3
30175 terrorismen 2
30176 terroristattack 2
30177 terroristbomber 1
30178 terrorister 6
30179 terroristerna 2
30180 terroristhandlingar 1
30181 terrorstyrka 1
30182 terräng 2
30183 terrängen 2
30184 tesen 2
30185 teservis 1
30186 testa 2
30187 testcentrer 1
30188 tester 1
30189 testet 1
30190 teve 1
30191 text 50
30192 texten 50
30193 textens 1
30194 texter 11
30195 texterna 5
30196 texternas 1
30197 textilsektorn 1
30198 textredigerare 2
30199 textändring 1
30200 that 1
30201 thatcherianska 1
30202 the 26
30203 therefore 1
30204 tibetaner 1
30205 tibetanerna 3
30206 tibetanska 5
30207 tid 212
30208 tiden 142
30209 tidens 6
30210 tider 14
30211 tiderna 1
30212 tidevarv 2
30213 tidig 5
30214 tidiga 9
30215 tidigare 222
30216 tidigarelagda 1
30217 tidigareläggas 1
30218 tidigt 23
30219 tidlöshet 1
30220 tidning 3
30221 tidningar 4
30222 tidningarna 2
30223 tidningen 5
30224 tidningsartikel 2
30225 tidplanen 1
30226 tidpunkt 21
30227 tidpunkten 9
30228 tidpunkter 1
30229 tids 4
30230 tidsaspekt 1
30231 tidsbegränsade 1
30232 tidsbegränsningen 3
30233 tidsbestämda 2
30234 tidsbestämmas 1
30235 tidsbrist 2
30236 tidsfaktorn 1
30237 tidsfrist 10
30238 tidsfristen 6
30239 tidsfristens 1
30240 tidsfrister 9
30241 tidsglappet 1
30242 tidsgräns 1
30243 tidshorisont 1
30244 tidsinställd 2
30245 tidsmässiga 2
30246 tidsperiod 6
30247 tidsperioder 1
30248 tidsplan 9
30249 tidsplanen 7
30250 tidspress 1
30251 tidsproblematiken 1
30252 tidsram 1
30253 tidsramar 5
30254 tidsramarna 2
30255 tidsramen 1
30256 tidsrymd 3
30257 tidsrymden 1
30258 tidsschemat 2
30259 tidsskede 1
30260 tidsskäl 1
30261 tidsskänken 1
30262 tidsålder 2
30263 tidsåtgång 1
30264 tidsödande 1
30265 tidtabell 17
30266 tidtabellen 2
30267 tidvatten 3
30268 tidvattnet 1
30269 tiga 2
30270 tigande 1
30271 tiger 5
30272 tigern 1
30273 tiggde 1
30274 tigger 1
30275 till 5961
30276 tillade 3
30277 tillbad 1
30278 tillbaka 168
30279 tillbakablick 1
30280 tillbakadragande 2
30281 tillbakadragandet 2
30282 tillbakadragen 1
30283 tillbakadragna 1
30284 tillbakagång 13
30285 tillbakalutad 1
30286 tillbakavisa 3
30287 tillbakavisande 2
30288 tillbakavisar 5
30289 tillbakavisat 1
30290 tillbakavisats 2
30291 tillbaks 4
30292 tillbehör 1
30293 tillblivelse 1
30294 tillbringa 3
30295 tillbringade 1
30296 tillbringat 3
30297 tillbud 1
30298 tillbörligt 1
30299 tilldela 2
30300 tilldelad 1
30301 tilldelade 1
30302 tilldelades 4
30303 tilldelar 2
30304 tilldelas 7
30305 tilldelats 7
30306 tilldelning 5
30307 tilldelningen 2
30308 tilldragelse 1
30309 tillerkände 1
30310 tillerkänner 3
30311 tillerkänns 1
30312 tillfalla 1
30313 tillfaller 1
30314 tillfinnandes 1
30315 tillflyktsort 1
30316 tillfoga 7
30317 tillfogar 1
30318 tillfogat 1
30319 tillfogats 1
30320 tillfreds 3
30321 tillfredsställa 4
30322 tillfredsställande 29
30323 tillfredsställde 1
30324 tillfredsställelse 13
30325 tillfrågats 1
30326 tillfälle 67
30327 tillfällen 41
30328 tillfället 32
30329 tillfällig 7
30330 tillfälliga 8
30331 tillfällighet 11
30332 tillfälligheter 1
30333 tillfälligt 12
30334 tillfälligtvis 1
30335 tillfångatagande 1
30336 tillför 9
30337 tillföra 8
30338 tillföras 1
30339 tillförlitlig 3
30340 tillförlitliga 4
30341 tillförlitlighet 2
30342 tillförlitlighetsproblem 1
30343 tillförlitligt 2
30344 tillförordnad 2
30345 tillförs 1
30346 tillförsikt 5
30347 tillförsäkra 1
30348 tillförsäkrar 1
30349 tillfört 1
30350 tillgivenhet 4
30351 tillgivet 1
30352 tillgodoräkna 1
30353 tillgodose 4
30354 tillgodosedda 2
30355 tillgodoser 1
30356 tillgodoses 3
30357 tillgripa 3
30358 tillgripas 1
30359 tillgriper 2
30360 tillgänglig 15
30361 tillgängliga 45
30362 tillgänglighet 3
30363 tillgängligheten 3
30364 tillgängligt 8
30365 tillgå 2
30366 tillgång 76
30367 tillgångar 10
30368 tillgången 18
30369 tillhandahålla 32
30370 tillhandahållande 25
30371 tillhandahållandet 2
30372 tillhandahållas 5
30373 tillhandahåller 12
30374 tillhandahållit 2
30375 tillhandahållits 5
30376 tillhandahållna 1
30377 tillhandahålls 3
30378 tillhandahöll 2
30379 tillhåll 1
30380 tillhör 31
30381 tillhöra 6
30382 tillhörande 2
30383 tillhörde 5
30384 tillhörighet 2
30385 tillhörigheten 2
30386 tillhörigheter 2
30387 tillika 3
30388 tillintetgjorts 1
30389 tillintetgöra 1
30390 tillit 2
30391 tillkom 3
30392 tillkommande 1
30393 tillkommer 9
30394 tillkommit 5
30395 tillkomst 2
30396 tillkomsten 1
30397 tillkrånglade 1
30398 tillkännagav 4
30399 tillkännage 2
30400 tillkännager 7
30401 tillkännages 3
30402 tillkännagett 1
30403 tillkännagivanden 3
30404 tillkännagivandena 1
30405 tillkännagivit 2
30406 tillkännagivits 1
30407 tillkännagivna 1
30408 tillmätas 1
30409 tillmäter 2
30410 tillmäts 2
30411 tillmötes 1
30412 tillmötesgå 2
30413 tillmötesgående 3
30414 tillmötesgås 1
30415 tillmötesgått 1
30416 tillnärmelsevis 1
30417 tillnärmning 11
30418 tillnärmningen 1
30419 tillnärmningsprocess 1
30420 tillrop 1
30421 tillryggalagt 1
30422 tillryggalagts 1
30423 tillryggalägger 1
30424 tillräcklig 39
30425 tillräckliga 17
30426 tillräckligt 110
30427 tillrätta 2
30428 tillrättalägger 1
30429 tillrättavisare 1
30430 tillrådligt 1
30431 tills 30
30432 tillsammans 150
30433 tillsats 3
30434 tillsatsdirektivet 1
30435 tillsatser 18
30436 tillsatserna 3
30437 tillsatsernas 1
30438 tillsatsämnen 1
30439 tillsatt 2
30440 tillsattes 1
30441 tillsatts 1
30442 tillse 13
30443 tillskansa 2
30444 tillskansar 1
30445 tillskapade 1
30446 tillskapandet 1
30447 tillskott 6
30448 tillskriver 2
30449 tillskrivs 1
30450 tillskyndar 2
30451 tillsluta 1
30452 tillstymmelse 1
30453 tillställa 1
30454 tillställningar 1
30455 tillställningarna 2
30456 tillställningen 2
30457 tillstå 2
30458 tillstånd 34
30459 tillstånden 2
30460 tillståndet 8
30461 tillståndsförfarandena 1
30462 tillståndssystem 1
30463 tillstår 1
30464 tillstås 1
30465 tillsyn 4
30466 tillsynsmyndighetens 1
30467 tillsynsmyndigheter 1
30468 tillsätt 1
30469 tillsätta 3
30470 tillsättandet 2
30471 tillsätter 1
30472 tillsättning 1
30473 tillsättningar 1
30474 tillsätts 3
30475 tillta 1
30476 tilltagande 2
30477 tilltal 1
30478 tilltala 1
30479 tilltalade 2
30480 tilltalande 1
30481 tilltalar 3
30482 tilltar 1
30483 tilltro 2
30484 tilltron 1
30485 tillträdandet 1
30486 tillträdde 1
30487 tillträde 29
30488 tillträdet 4
30489 tilltänkta 1
30490 tillval 1
30491 tillvara 3
30492 tillvarata 1
30493 tillvaro 8
30494 tillvaron 2
30495 tillverka 5
30496 tillverkade 1
30497 tillverkar 3
30498 tillverkaransvar 1
30499 tillverkaransvaret 4
30500 tillverkare 3
30501 tillverkaren 11
30502 tillverkarens 2
30503 tillverkarna 15
30504 tillverkarnas 6
30505 tillverkas 4
30506 tillverkats 2
30507 tillverkning 3
30508 tillverkningen 4
30509 tillverkningsindustri 1
30510 tillverkningsindustrin 5
30511 tillverkningsprocesser 1
30512 tillverkningssektorn 2
30513 tillväga 6
30514 tillvägagångssätt 23
30515 tillvägagångssätten 1
30516 tillvägagångssättet 4
30517 tillväxt 77
30518 tillväxt- 2
30519 tillväxtbefrämjande 1
30520 tillväxtbranscherna 1
30521 tillväxtcentrum 1
30522 tillväxtdynamik 1
30523 tillväxten 30
30524 tillväxtfaktor 1
30525 tillväxtfaktorer 1
30526 tillväxtmål 2
30527 tillväxtmålsättningar 1
30528 tillväxtnivå 4
30529 tillväxtnivåer 1
30530 tillväxtpotential 1
30531 tillväxtprognosen 1
30532 tillväxttakt 2
30533 tillväxtökande 1
30534 tillägg 15
30535 tillägga 21
30536 tillägget 1
30537 tilläggs 1
30538 tilläggsbudget 1
30539 tilläggsfråga 3
30540 tilläggskrav 1
30541 tillägna 2
30542 tillämpa 82
30543 tillämpad 1
30544 tillämpades 1
30545 tillämpande 1
30546 tillämpandet 1
30547 tillämpar 16
30548 tillämpas 91
30549 tillämpat 2
30550 tillämpats 9
30551 tillämplig 7
30552 tillämpliga 9
30553 tillämplighet 2
30554 tillämpligt 4
30555 tillämpning 63
30556 tillämpningar 1
30557 tillämpningarna 1
30558 tillämpningen 61
30559 tillämpningsbestämmelser 1
30560 tillämpningsbestämmelserna 2
30561 tillämpningsförfaranden 1
30562 tillämpningsförordning 1
30563 tillämpningsförordningen 2
30564 tillämpningsområde 6
30565 tillämpningsområdet 6
30566 tillämpningsprocessen 1
30567 tillämpningsstrategier 1
30568 tillämpningssvårigheter 1
30569 tillämpningsövervakning 1
30570 tillät 1
30571 tillåt 2
30572 tillåta 35
30573 tillåtande 1
30574 tillåtas 13
30575 tillåtelse 1
30576 tillåten 6
30577 tillåter 49
30578 tillåtet 4
30579 tillåtits 1
30580 tillåtliga 1
30581 tillåtna 12
30582 tillåts 11
30583 timing 1
30584 timjan 1
30585 timma 1
30586 timmar 27
30587 timmarna 1
30588 timmars 1
30589 timme 14
30590 ting 19
30591 tingens 1
30592 tinninglockar 2
30593 tinningådror 1
30594 tio 54
30595 tionde 1
30596 tionyheterna 1
30597 tiopundssedlarna 1
30598 tiotal 3
30599 tiotals 8
30600 tiotusen 1
30601 tiotusentals 5
30602 tioårsperioden 1
30603 tips 2
30604 tisdag 2
30605 tisdagen 2
30606 tisdagens 1
30607 titan 1
30608 titel 2
30609 titeln 10
30610 titelsektionen 1
30611 titlar 1
30612 titt 6
30613 titta 53
30614 tittade 20
30615 tittande 2
30616 tittar 20
30617 tittarnöje 1
30618 tja 1
30619 tjata 1
30620 tjatig 1
30621 tjeckiske 2
30622 tjejer 1
30623 tjetjenska 4
30624 tjetjenskt 2
30625 tjock 4
30626 tjocka 5
30627 tjockisen 1
30628 tjockleken 1
30629 tjockolja 2
30630 tjugo 10
30631 tjugofem 5
30632 tjugoförsta 2
30633 tjugonde 4
30634 tjugosex 1
30635 tjugosexåriga 1
30636 tjugosju 2
30637 tjugotusen 2
30638 tjugotvå 1
30639 tjugotvåtusen 1
30640 tjugu 1
30641 tjur 1
30642 tjuren 2
30643 tjurskallig 1
30644 tjusade 1
30645 tjusar 1
30646 tjusat 1
30647 tjusig 2
30648 tjusning 1
30649 tjuvnad 1
30650 tjäna 14
30651 tjänade 1
30652 tjänar 26
30653 tjänare 1
30654 tjänaren 1
30655 tjänarstaben 1
30656 tjänas 1
30657 tjänat 5
30658 tjänst 35
30659 tjänstberett 1
30660 tjänsteenhet 1
30661 tjänsteenheter 4
30662 tjänsteenheterna 1
30663 tjänstefel 1
30664 tjänsteföreskrifterna 6
30665 tjänsteföretag 1
30666 tjänsteföretagen 2
30667 tjänstekriterier 1
30668 tjänstekvaliteten 3
30669 tjänsteleverantören 2
30670 tjänsteman 9
30671 tjänstemanna-apparaten 1
30672 tjänstemannakårer 1
30673 tjänstemannarepresentanter 1
30674 tjänstemän 42
30675 tjänstemännen 11
30676 tjänstemännens 4
30677 tjänstemäns 3
30678 tjänsten 6
30679 tjänstenivå 5
30680 tjänstenivån 2
30681 tjänstens 1
30682 tjänsteproducenter 3
30683 tjänsteproducenterna 1
30684 tjänsteproducenters 1
30685 tjänsteproduktion 1
30686 tjänster 109
30687 tjänsterna 22
30688 tjänsternas 1
30689 tjänsterum 1
30690 tjänstesektorer 1
30691 tjänstesektorn 4
30692 tjänsteuppdrag 2
30693 tjänsteutbudet 1
30694 tjänsteåligganden 1
30695 tjänstgjorde 1
30696 tjänstgjort 1
30697 tjänstgör 1
30698 tjänstgörande 15
30699 tjära 2
30700 tjöt 1
30701 to 2
30702 toalettbord 1
30703 toaletten 2
30704 toaletter 1
30705 toaletterna 2
30706 toalettköerna 1
30707 tobak 1
30708 tobaksblommorna 1
30709 tobaksodling 1
30710 tobakspung 1
30711 toddyn 1
30712 todo 1
30713 tofflorna 1
30714 tofsar 1
30715 tog 115
30716 toga 1
30717 togorna 1
30718 togs 23
30719 tokig 2
30720 tolerans 15
30721 toleransen 1
30722 toleranskulturen 1
30723 tolerant 1
30724 toleranta 3
30725 tolerera 3
30726 tolererar 1
30727 tolereras 7
30728 tolk 1
30729 tolka 8
30730 tolkade 3
30731 tolkar 10
30732 tolkarna 4
30733 tolkarnas 1
30734 tolkas 13
30735 tolkat 1
30736 tolkats 2
30737 tolkning 20
30738 tolkningar 4
30739 tolkningarna 1
30740 tolkningarnas 1
30741 tolkningen 10
30742 tolkningsmeddelanden 1
30743 tolkningsmöjligheterna 1
30744 tolkningsproblem 1
30745 tolv 6
30746 tom 5
30747 tomater 3
30748 tomatkonserver 1
30749 tomatpuré 1
30750 tomhet 3
30751 tomma 7
30752 tomrum 5
30753 ton 34
30754 toner 1
30755 tonfall 4
30756 tonfisk 18
30757 tonfiskbestånden 1
30758 tonfisken 5
30759 tonfisket 1
30760 tonfiskliknande 1
30761 tongivande 1
30762 tongångar 1
30763 tonlös 1
30764 tonvikt 6
30765 tonvikten 3
30766 tonåringar 1
30767 tonårsgrammofonen 1
30768 topp 3
30769 toppen 7
30770 toppluva 1
30771 toppmöte 14
30772 toppmöten 3
30773 toppmötena 1
30774 toppmötesnivå 1
30775 toppmötet 73
30776 toppnyhet 1
30777 toppositioner 1
30778 topprioritet 1
30779 topptjänstemän 1
30780 torde 5
30781 tordönsröst 1
30782 torftig 1
30783 torg 1
30784 torka 12
30785 torkade 3
30786 torkan 1
30787 torkas 1
30788 torkat 1
30789 torna 1
30790 tornet 1
30791 torniga 1
30792 torpet 2
30793 torra 4
30794 torrare 1
30795 torrlägger 1
30796 torrt 1
30797 torsdag 15
30798 torsdagen 7
30799 torsdagens 1
30800 torsdags 1
30801 torsk 3
30802 torskbestånden 1
30803 torsken 1
30804 torskfiske 1
30805 torskkvot 1
30806 torskkvoten 1
30807 torteras 2
30808 torterats 1
30809 tortyr 4
30810 tortyren 1
30811 tortyrinstrument 1
30812 torven 4
30813 torvvatten 1
30814 total 13
30815 totala 35
30816 totalanslag 2
30817 totalanslaget 3
30818 totalansvar 1
30819 totalbeloppet 1
30820 totalblockad 1
30821 totalfångst 2
30822 totalfångsten 2
30823 totalförbud 2
30824 totalförstört 1
30825 totalitarism 2
30826 totalitarismens 1
30827 totalitära 2
30828 totalsumma 1
30829 totalsumman 1
30830 totalt 22
30831 totalvolym 1
30832 toxiska 1
30833 trader 1
30834 tradition 15
30835 traditionalism 1
30836 traditionell 4
30837 traditionella 16
30838 traditionellt 4
30839 traditionen 5
30840 traditionens 1
30841 traditioner 8
30842 traditionerna 2
30843 trafik 5
30844 trafik- 1
30845 trafikanter 1
30846 trafikeländet 1
30847 trafiken 7
30848 trafikens 1
30849 trafikerar 1
30850 trafikkontroller 1
30851 trafikled 1
30852 trafikolyckor 1
30853 trafikpolisen 1
30854 trafikpoliser 1
30855 trafikstockningar 1
30856 trafiksäkerhet 1
30857 trafiksäkerheten 8
30858 tragedi 10
30859 tragedier 6
30860 tragedin 6
30861 tragisk 3
30862 tragiska 12
30863 tragiskt 8
30864 trakasserier 3
30865 trakt 1
30866 trakten 1
30867 trakterna 1
30868 tramp 1
30869 trampar 1
30870 trans 3
30871 transaktioner 2
30872 transaktionskostnader 1
30873 transatlantiska 2
30874 transeuropeiska 7
30875 transferable 2
30876 transfereringar 1
30877 transformera 2
30878 transformeras 3
30879 transithallen 1
30880 transitivt 1
30881 transitland 2
30882 transitländer 1
30883 transitrutten 1
30884 transittrafiken 1
30885 transmissibel 1
30886 transnationell 3
30887 transnationella 6
30888 transnationellt 4
30889 transport 78
30890 transport- 5
30891 transportabla 1
30892 transportbeställarna 1
30893 transportbestämmelser 1
30894 transportdirektiv 1
30895 transporten 7
30896 transporter 27
30897 transportera 3
30898 transporterade 2
30899 transporterades 1
30900 transporterar 2
30901 transporteras 8
30902 transporterna 5
30903 transportfederationen 1
30904 transportfrågor 1
30905 transportgruppen 1
30906 transportkapacitet 1
30907 transportkostnaderna 2
30908 transportmarknad 1
30909 transportmedel 1
30910 transportministrar 1
30911 transportnät 3
30912 transportnäten 2
30913 transportområden 1
30914 transportområdet 2
30915 transportpolitik 1
30916 transportpolitiken 2
30917 transportpolitiker 1
30918 transportpolitiska 1
30919 transportproblem 1
30920 transportsektorn 2
30921 transportsäkerhet 3
30922 transportsäkerheten 3
30923 transportsätt 1
30924 transportutskottet 1
30925 transportörernas 1
30926 trappa 1
30927 trappan 10
30928 trappavsatsen 2
30929 trapphallen 1
30930 trappsteg 1
30931 trappsteget 1
30932 trasa 1
30933 trasas 1
30934 trasig 2
30935 trasiga 4
30936 trasigt 1
30937 trasmatta 1
30938 trasmattan 1
30939 trasor 1
30940 trassel 1
30941 trassla 1
30942 trasslade 2
30943 trasslat 1
30944 trasslig 1
30945 traumatiska 1
30946 travar 3
30947 traven 2
30948 travesterade 1
30949 tre 172
30950 tre-fyra 1
30951 trea 1
30952 trebent 1
30953 tredagarskryssning 1
30954 tredelade 1
30955 tredje 187
30956 tredjedel 12
30957 tredjedelar 4
30958 tredjelandsmedborgare 6
30959 tredjelandsmedborgares 1
30960 trehjulingar 1
30961 trehundrafemti 1
30962 trekilometerspromenad 1
30963 treklang 1
30964 tremånadersfristen 1
30965 tremånadersperioden 2
30966 trend 4
30967 trenden 3
30968 trender 1
30969 trepartsagerande 1
30970 trepartsarbete 1
30971 trepartsarbetsgrupp 3
30972 trepartsarbetsgruppen 1
30973 trepartsmöte 1
30974 trepartssamtalen 1
30975 trephena-mat 1
30976 treprocentsnormen 1
30977 trettio 12
30978 trettiofem 3
30979 trettiofemårsåldern 1
30980 trettiotal 1
30981 trettiotalet 3
30982 trettioåtta 1
30983 tretton 6
30984 trettonde 1
30985 trettonåriga 1
30986 trevlig 2
30987 trevligt 5
30988 treårsperioder 1
30989 triangel 1
30990 triangelformad 1
30991 triangelförhållande 1
30992 tribunal 2
30993 tribunen 1
30994 tributyl 1
30995 trick 1
30996 trikåfabrik 1
30997 trilbyhatt 1
30998 triljoner 1
30999 trimmade 1
31000 trio 1
31001 trirem 1
31002 trist 5
31003 trista 1
31004 triumf 1
31005 triumferat 1
31006 trivas 1
31007 trivdes 3
31008 trivialaste 1
31009 trivsamma 1
31010 tro 62
31011 trodde 20
31012 trofasthet 1
31013 troféer 1
31014 trogen 5
31015 troget 2
31016 trogne 1
31017 trojanska 1
31018 trojkan 1
31019 troliga 1
31020 troligen 10
31021 troligt 6
31022 troligtvis 4
31023 trolldom 1
31024 trolldomsböcker 1
31025 trolldomskraft 1
31026 trolleri 1
31027 trolleriet 1
31028 trollguld 1
31029 trollkarl 4
31030 trollkarlar 3
31031 trollkarlsbutik 1
31032 trollkarlshatt 1
31033 trollkarlshem 1
31034 trollkarlsskolan 1
31035 trollkarlsvärlden 3
31036 trollkonst 1
31037 trollspö 2
31038 trollspöt 1
31039 trollstav 3
31040 trollstaven 1
31041 tron 1
31042 tropisk 1
31043 tropiska 15
31044 tror 485
31045 trosartikel 1
31046 trots 152
31047 trott 7
31048 trottoaren 2
31049 trottoarer 1
31050 trottoarerna 1
31051 trovärdig 8
31052 trovärdiga 8
31053 trovärdige 1
31054 trovärdighet 29
31055 trovärdigheten 4
31056 trovärdighetskris 1
31057 trovärdighetsproblem 1
31058 trovärdighetstest 1
31059 trovärdighetstestet 1
31060 trovärdigt 2
31061 trubbigt 1
31062 trumfkort 3
31063 trummade 1
31064 trumpet 1
31065 trumpinnar 1
31066 trupper 8
31067 truppminor 1
31068 trusten 1
31069 truster 2
31070 trusterna 1
31071 tryck 14
31072 trycka 6
31073 tryckalster 1
31074 tryckas 1
31075 tryckbärande 1
31076 trycker 2
31077 trycket 8
31078 tryckfel 1
31079 tryckfriheten 1
31080 tryckningen 1
31081 tryckta 2
31082 tryckte 6
31083 trygg 1
31084 trygga 3
31085 tryggad 1
31086 tryggande 1
31087 tryggas 1
31088 trygghet 52
31089 tryggheten 37
31090 trygghetsmodellen 1
31091 trygghetsnivå 1
31092 trygghetspolitik 1
31093 trygghetssystem 9
31094 trygghetssystemen 21
31095 trygghetssystemens 3
31096 trygghetssystemet 4
31097 tryggt 3
31098 trä 4
31099 träbord 1
31100 träd 10
31101 träda 19
31102 trädde 13
31103 träddungar 1
31104 träddunge 1
31105 träden 5
31106 träder 12
31107 trädgårdar 2
31108 trädgården 5
31109 trädgårdsanläggningarna 1
31110 trädgårdsbänken 3
31111 trädgårdshäcken 1
31112 trädgårdsmöbeln 1
31113 trädgårdsprodukter 1
31114 trädgårdsstolarna 1
31115 trädstruktur 1
31116 trädtopparna 1
31117 träffa 13
31118 träffade 13
31119 träffades 4
31120 träffande 3
31121 träffar 7
31122 träffas 8
31123 träffat 2
31124 träffats 2
31125 träkolsgrill 1
31126 träldom 2
31127 trälåda 1
31128 tränat 1
31129 tränga 2
31130 trängande 1
31131 trängde 5
31132 trängdes 1
31133 tränger 4
31134 trängt 2
31135 träning 1
31136 träproduktion 1
31137 träsk 2
31138 träskulpturerna 1
31139 träskylt 1
31140 trätor 1
31141 trätt 10
31142 tråd 3
31143 trådar 4
31144 trådarna 1
31145 trådde 1
31146 tråden 2
31147 tråkigaste 1
31148 tråkigt 8
31149 trålar 1
31150 trånga 1
31151 trångmål 1
31152 trångt 1
31153 tröga 2
31154 tröghet 5
31155 trögheten 2
31156 tröskade 1
31157 tröskel 3
31158 tröskeln 5
31159 tröskelvärdet 1
31160 tröst 3
31161 tröstad 1
31162 tröstade 1
31163 tröstegrund 1
31164 trött 6
31165 trötta 3
31166 trötthet 2
31167 tröttnade 2
31168 tröttsamma 1
31169 tröttsamt 1
31170 tsetseflugor 1
31171 tudelad 1
31172 tuff 1
31173 tuffare 1
31174 tuffingarna 1
31175 tufft 2
31176 tull 2
31177 tull- 1
31178 tullavgifter 1
31179 tullavgifterna 1
31180 tullförvaltningen 1
31181 tullgåvor 1
31182 tullhinder 1
31183 tullintegration 1
31184 tullkontroll 1
31185 tullmyndighet 1
31186 tullmyndigheten 1
31187 tullmyndigheter 1
31188 tullmyndigheterna 3
31189 tullsamarbetskommittén 1
31190 tulltariff 1
31191 tulltjänstemän 2
31192 tulltjänstemännen 1
31193 tulltjänstemännens 1
31194 tulltjänster 1
31195 tullättnader 1
31196 tumma 3
31197 tummarna 1
31198 tummen 1
31199 tumultet 1
31200 tumultuarisk 1
31201 tunc 1
31202 tung 15
31203 tunga 12
31204 tungmetaller 8
31205 tungmetallerna 1
31206 tungrodd 1
31207 tungrodda 1
31208 tungroddhet 1
31209 tungsint 1
31210 tungt 8
31211 tunna 3
31212 tunnades 1
31213 tunneln 2
31214 tunneltrafik 1
31215 tunnland 2
31216 tunnlar 2
31217 tunnlarna 1
31218 tunt 3
31219 tur 29
31220 turer 1
31221 turism 70
31222 turismen 50
31223 turismens 4
31224 turismfrågor 1
31225 turista 1
31226 turistbranschen 2
31227 turistbyråerna 1
31228 turistcentrer 2
31229 turister 4
31230 turisterna 2
31231 turisthandel 1
31232 turistindustri 1
31233 turistindustrin 6
31234 turistiskt 2
31235 turistland 1
31236 turistmarknaden 3
31237 turistmål 1
31238 turistmålet 1
31239 turistnäring 4
31240 turistnäringen 18
31241 turistnäringens 4
31242 turistområde 1
31243 turistområdet 1
31244 turistorterna 1
31245 turistpolitik 3
31246 turistpolitiken 2
31247 turistpotential 1
31248 turistsektorers 1
31249 turistsektorn 5
31250 turistsäsongen 2
31251 turistutbildningen 1
31252 turkar 2
31253 turkarna 2
31254 turkarnas 1
31255 turkcyprioter 1
31256 turkcyprioterna 1
31257 turkcypriotiska 6
31258 turkcypriotiske 1
31259 turkisk-grekiska 1
31260 turkiska 20
31261 turkiske 3
31262 turn-over 1
31263 tusan 2
31264 tusen 17
31265 tusentals 24
31266 tuta 1
31267 tutade 2
31268 tveka 5
31269 tvekade 1
31270 tvekan 42
31271 tvekar 8
31272 tvekat 2
31273 tveklöst 4
31274 tveksam 5
31275 tveksamhet 2
31276 tveksamma 2
31277 tveksamt 3
31278 tvetydig 3
31279 tvetydiga 3
31280 tvetydighet 5
31281 tvetydigheten 1
31282 tvetydigheter 1
31283 tvillingarna 1
31284 tvillingbröder 1
31285 tvillingpar 1
31286 tvinga 15
31287 tvingad 2
31288 tvingade 6
31289 tvingades 5
31290 tvingande 11
31291 tvingar 15
31292 tvingas 27
31293 tvingats 4
31294 tvinnade 2
31295 tvist 4
31296 tvista 1
31297 tvistefrågor 1
31298 tvisten 1
31299 tvister 6
31300 tvivel 66
31301 tvivelaktig 3
31302 tvivelaktiga 2
31303 tvivelsmålen 1
31304 tvivelsutan 3
31305 tvivla 1
31306 tvivlar 17
31307 tvivlat 1
31308 tvungen 28
31309 tvungna 22
31310 tvärgående 2
31311 tvärpolitiska 2
31312 tvärs 7
31313 tvärsöver 1
31314 tvärt 2
31315 tvärtemot 4
31316 tvärtom 36
31317 tvätta 3
31318 tvättade 2
31319 tvättat 1
31320 tvättfat 1
31321 tvättmedelseksem 1
31322 två 412
31323 två-ett 1
31324 två-tre 1
31325 tvåhundra 5
31326 tvåhundraåriga 1
31327 tvålbit 1
31328 tvålflingor 1
31329 tvång 5
31330 tvånget 3
31331 tvångsarbetarna 2
31332 tvångsfinansieras 1
31333 tvångsförflyttade 2
31334 tvångsförflyttats 2
31335 tvångsintegrerats 1
31336 tvångsmarschen 1
31337 tvångsmedel 1
31338 tvångsmekanism 1
31339 tvångsrekryteras 1
31340 tvångsstruktur 1
31341 tvångströja 1
31342 tvångströjor 1
31343 tvåprocentströskeln 1
31344 tvåspråksutbildningen 1
31345 tvåtusen 1
31346 tvåårig 1
31347 tvååriga 1
31348 twist 1
31349 ty 31
31350 tycka 6
31351 tyckas 3
31352 tycke 4
31353 tycker 196
31354 tycks 32
31355 tyckt 5
31356 tyckte 25
31357 tycktes 18
31358 tyckts 1
31359 tydde 1
31360 tyder 13
31361 tydlig 44
31362 tydliga 44
31363 tydligare 19
31364 tydligaste 3
31365 tydligen 15
31366 tydliggjorde 1
31367 tydliggjort 2
31368 tydliggör 4
31369 tydliggöra 4
31370 tydliggöras 1
31371 tydliggörs 1
31372 tydlighet 10
31373 tydligt 166
31374 tyg 1
31375 tygellösa 1
31376 tygla 1
31377 tygleksaker 1
31378 tynande 1
31379 tynga 2
31380 tyngande 1
31381 tyngas 1
31382 tyngd 7
31383 tyngdpunkt 1
31384 tyngdpunkten 3
31385 tyngdpunkter 1
31386 tynger 3
31387 tyngre 1
31388 tyngst 1
31389 tyngsta 1
31390 typ 70
31391 typen 36
31392 typer 19
31393 typerna 2
31394 typexempel 1
31395 typfall 1
31396 typgodkännanden 1
31397 typiska 1
31398 typiskt 2
31399 typtrogen 1
31400 tyranners 1
31401 tyranni 4
31402 tysk 2
31403 tyska 33
31404 tyskar 1
31405 tyskarna 1
31406 tyske 3
31407 tyskspråkig 1
31408 tyskt 2
31409 tyst 16
31410 tysta 6
31411 tystar 1
31412 tystare 2
31413 tystlåten 1
31414 tystnad 12
31415 tystnade 3
31416 tystnaden 1
31417 tystnar 1
31418 tyvärr 79
31419 täcka 6
31420 täckande 1
31421 täckas 2
31422 täcker 18
31423 täckmantel 1
31424 täcks 8
31425 täckt 1
31426 täckte 1
31427 tält 2
31428 tältet 2
31429 tämligen 7
31430 tända 1
31431 tändanordningarna 1
31432 tändas 1
31433 tände 3
31434 tänder 4
31435 tänderna 1
31436 tändes 2
31437 tänds 1
31438 tändsticka 1
31439 tändstickor 2
31440 tänja 1
31441 tänjas 1
31442 tänk 6
31443 tänka 89
31444 tänkande 1
31445 tänkandet 2
31446 tänkas 8
31447 tänkbar 1
31448 tänkbara 9
31449 tänkbart 2
31450 tänker 113
31451 tänkesättet 1
31452 tänkt 15
31453 tänkta 2
31454 tänkte 26
31455 tänktes 1
31456 tänkvärt 1
31457 tänt 1
31458 täppa 4
31459 täpper 1
31460 tärningsspel 1
31461 tärt 2
31462 täta 3
31463 tätare 2
31464 tätbefolkat 2
31465 täten 3
31466 tätortsområden 1
31467 tätt 3
31468 tävla 1
31469 tävlade 1
31470 tävlar 2
31471 tävling 2
31472 tå 4
31473 tåg 5
31474 tåg- 1
31475 tåget 3
31476 tågets 1
31477 tågkraschen 1
31478 tågolyckan 1
31479 tål 1
31480 tålamod 4
31481 tålig 1
31482 tåligt 1
31483 tålmodigt 1
31484 tårstrimmiga 1
31485 tårta 2
31486 töckniga 1
31487 töcknigt 1
31488 tömd 1
31489 tömma 1
31490 tömmer 1
31491 töms 4
31492 tömt 1
31493 törs 1
31494 u-länderna 4
31495 u-ländernas 1
31496 udda 2
31497 uggla 3
31498 ugglan 1
31499 ugglor 1
31500 ugnen 1
31501 ultimatum 1
31502 ultraliberala 4
31503 ultraliberalism 1
31504 ultraperifer 1
31505 ultraperifera 2
31506 umbärande 1
31507 umgänge 1
31508 umgängesformer 1
31509 umgänget 1
31510 umgåtts 1
31511 un 2
31512 una 2
31513 und 1
31514 undan 26
31515 undanber 2
31516 undandrar 1
31517 undandras 1
31518 undanflykter 2
31519 undanforslad 1
31520 undanglidande 1
31521 undanhålla 2
31522 undanmanövrar 1
31523 undanröja 12
31524 undanröjas 1
31525 undanröjer 1
31526 undanröjts 1
31527 undanslagna 1
31528 undanta 6
31529 undantag 59
31530 undantagen 6
31531 undantaget 6
31532 undantagna 3
31533 undantagsbestämmelser 1
31534 undantagsfall 2
31535 undantagsförfarandet 1
31536 undantagsförordning 1
31537 undantagsmässig 1
31538 undantagsperiod 1
31539 undantagsregeln 3
31540 undantagsregler 1
31541 undantagssituationer 1
31542 undantagstillstånd 1
31543 undantagstillståndet 1
31544 undantagsvis 1
31545 undantas 4
31546 under 893
31547 underarmen 1
31548 underbar 3
31549 underbara 1
31550 underbart 4
31551 underblåsa 1
31552 underblåser 3
31553 underbygga 1
31554 underbyggda 2
31555 undercover-verksamhet 1
31556 underfinansierade 1
31557 underformulär 1
31558 underfund 3
31559 underförstådd 1
31560 underförstås 1
31561 underförstått 1
31562 undergräva 5
31563 undergrävas 3
31564 undergräver 3
31565 undergrävs 1
31566 undergång 1
31567 undergår 1
31568 underhandsrapport 1
31569 underhus 1
31570 underhuset 4
31571 underhåll 5
31572 underhåller 1
31573 underhållet 2
31574 underhållna 1
31575 underhållningsbranschen 1
31576 underhålls 1
31577 underjordiska 4
31578 underkasta 4
31579 underkastad 1
31580 underkastas 2
31581 underkastat 1
31582 underkastelse 1
31583 underkastelsen 1
31584 underkategori 2
31585 underlag 8
31586 underlaget 1
31587 underleverantörer 4
31588 underleverantörsområdet 1
31589 underlig 1
31590 underliga 2
31591 underliggande 9
31592 underligt 2
31593 underläge 2
31594 underlägset 1
31595 underlägsna 3
31596 underläpp 1
31597 underlätta 37
31598 underlättar 10
31599 underlättats 1
31600 underlåtande 1
31601 underlåtenhet 3
31602 underlåtenheten 1
31603 underlåter 4
31604 underlåtit 2
31605 undermappar 1
31606 undermeningen 1
31607 underminera 2
31608 underminerar 1
31609 undermineras 1
31610 undermålig 1
31611 undermåliga 1
31612 undernärda 1
31613 underordnad 2
31614 underordnade 2
31615 underordnande 1
31616 underordnas 4
31617 underordnat 1
31618 underprivilegierade 1
31619 underprogram 1
31620 underpunkt 4
31621 underrapporter 2
31622 underrepresentation 3
31623 underrepresentationen 1
31624 underrepresenterade 5
31625 underrätta 1
31626 underrättas 1
31627 underrättat 1
31628 underrättelsetjänst 1
31629 underrättelsetjänsten 1
31630 underrättelsetjänster 1
31631 underrättelsetjänsternas 1
31632 underrättelseverksamheten 1
31633 underskatta 2
31634 underskattad 1
31635 underskattade 1
31636 underskattas 2
31637 underskattat 1
31638 underskott 21
31639 underskotten 6
31640 underskottet 16
31641 underskrider 1
31642 underskrift 2
31643 underskrifter 1
31644 understiger 1
31645 understrukit 3
31646 understrukits 2
31647 understrukna 1
31648 understryka 46
31649 understrykas 5
31650 understryker 11
31651 understryks 7
31652 underströk 7
31653 underströks 1
31654 underström 1
31655 underställa 1
31656 underställas 4
31657 underställd 3
31658 underställda 2
31659 underställs 2
31660 underställt 2
31661 underställts 1
31662 understå 1
31663 understöd 1
31664 understöddes 1
31665 understöder 2
31666 understödja 3
31667 understödjande 1
31668 understödjas 3
31669 understöds 1
31670 understödspolitik 1
31671 undersysselsättningens 1
31672 undersåte 1
31673 undersöka 33
31674 undersökande 2
31675 undersökas 10
31676 undersöker 4
31677 undersökning 22
31678 undersökningar 20
31679 undersökningarna 3
31680 undersökningarnas 1
31681 undersökningen 7
31682 undersökningsgrupp 1
31683 undersökningskommission 1
31684 undersökningskommitté 1
31685 undersökningskommittén 1
31686 undersökningsmakt 1
31687 undersökningsmekanismer 1
31688 undersökningsprocess 2
31689 undersökningssystem 1
31690 undersökt 6
31691 undersökta 2
31692 undersökte 1
31693 underteckna 6
31694 undertecknad 1
31695 undertecknade 2
31696 undertecknades 9
31697 undertecknande 1
31698 undertecknandet 1
31699 undertecknar 5
31700 undertecknarna 1
31701 undertecknas 3
31702 undertecknat 17
31703 undertecknats 4
31704 undertrycka 3
31705 undertrycker 2
31706 undertryckta 1
31707 underutnyttjande 1
31708 underutvecklad 3
31709 underutvecklade 3
31710 underutvecklat 1
31711 underutveckling 2
31712 underutvecklingen 2
31713 undervattensfloder 1
31714 undervattenssamling 1
31715 undervegetationen 1
31716 underverk 1
31717 undervisa 1
31718 undervisning 3
31719 undervisningen 2
31720 undervärdera 1
31721 undfallande 1
31722 undgick 1
31723 undgå 2
31724 undgår 3
31725 undgått 3
31726 undkomma 2
31727 undkommer 2
31728 undkommit 2
31729 undlåtit 1
31730 undra 5
31731 undrade 9
31732 undran 4
31733 undrande 2
31734 undrar 39
31735 undsluppit 1
31736 undsätta 1
31737 undvik 1
31738 undvika 86
31739 undvikas 8
31740 undviker 8
31741 undvikit 4
31742 undvikits 1
31743 undviks 2
31744 ung 17
31745 ung. 1
31746 unga 35
31747 ungdom 3
31748 ungdomar 22
31749 ungdomarna 3
31750 ungdomarnas 1
31751 ungdomen 2
31752 ungdomlig 1
31753 ungdoms- 3
31754 ungdomsarbetslöshet 2
31755 ungdomsarbetslösheten 1
31756 ungdomsbrottslighet 3
31757 ungdomsfrågor 3
31758 unge 11
31759 ungefär 19
31760 ungefärliga 1
31761 ungerska 1
31762 ungfisken 1
31763 ungrare 1
31764 ungt 1
31765 uniform 2
31766 uniformer 1
31767 uniformerade 1
31768 unik 3
31769 unika 12
31770 unikt 6
31771 unilaterala 2
31772 unilateralt 3
31773 union 60
31774 unionen 854
31775 unionen-Afrika 2
31776 unionen-Kina 1
31777 unionens 406
31778 unions 1
31779 unions- 1
31780 unionsfördrag 1
31781 unionsfördraget 1
31782 unionsmedborgare 2
31783 unionsmedborgarna 1
31784 unionsmedborgarnas 2
31785 unionsmedlemmar 1
31786 unionsnivå 6
31787 unionssammanhang 1
31788 universalitet 1
31789 universaliteten 1
31790 universalmedel 1
31791 universell 3
31792 universella 10
31793 universitet 2
31794 universiteten 1
31795 universitetet 4
31796 universitetsmiljöerna 1
31797 universum 1
31798 universums 2
31799 unna 1
31800 uns 1
31801 unset 1
31802 upp 794
31803 uppassade 1
31804 uppassare 1
31805 uppbackning 1
31806 uppbjuda 1
31807 uppblandad 1
31808 uppblandning 1
31809 uppblötta 1
31810 uppborstat 1
31811 uppbringa 1
31812 uppbringar 2
31813 uppbringas 2
31814 uppbromsningen 1
31815 uppbrottsstämning 1
31816 uppburits 1
31817 uppbyggande 1
31818 uppbyggandet 1
31819 uppbyggd 1
31820 uppbyggnad 5
31821 uppbyggnaden 16
31822 uppbyggnadsplatserna 1
31823 uppbyggt 4
31824 uppbär 1
31825 uppbära 2
31826 uppbåda 2
31827 uppdatera 6
31828 uppdaterad 1
31829 uppdateras 1
31830 uppdatering 1
31831 uppdelade 1
31832 uppdelat 4
31833 uppdelning 4
31834 uppdelningen 3
31835 uppdrag 41
31836 uppdragen 1
31837 uppdraget 5
31838 uppdragna 1
31839 uppdrog 1
31840 uppdykandet 1
31841 uppe 16
31842 uppehälle 2
31843 uppehåll 2
31844 uppehålla 12
31845 uppehåller 4
31846 uppehållet 1
31847 uppehållit 1
31848 uppehållstillstånd 5
31849 uppehållstillståndet 2
31850 uppehållstillståndets 1
31851 uppehållsvillkor 1
31852 uppenbar 6
31853 uppenbara 6
31854 uppenbarar 1
31855 uppenbarelse 2
31856 uppenbarligen 29
31857 uppenbart 69
31858 uppfanns 1
31859 uppfatta 2
31860 uppfattade 4
31861 uppfattar 20
31862 uppfattas 6
31863 uppfattat 3
31864 uppfattbart 1
31865 uppfattning 71
31866 uppfattningar 10
31867 uppfattningen 13
31868 uppfinna 3
31869 uppfinning 1
31870 uppfinningarnas 1
31871 uppfostrades 1
31872 uppfostran 2
31873 uppfriskande 1
31874 uppfylla 60
31875 uppfyllandet 6
31876 uppfyllas 11
31877 uppfylld 2
31878 uppfyllda 4
31879 uppfyllde 3
31880 uppfylldes 2
31881 uppfyller 36
31882 uppfylls 8
31883 uppfyllt 1
31884 uppfyllts 5
31885 uppfångade 1
31886 uppfödning 1
31887 uppföljas 1
31888 uppföljning 15
31889 uppföljningen 6
31890 uppföljningsfråga 1
31891 uppföljningskommittén 2
31892 uppföljningsrapporten 1
31893 uppföljningsregler 1
31894 uppför 11
31895 uppföra 4
31896 uppförande 5
31897 uppförandekod 6
31898 uppförandekoden 3
31899 uppförandekoder 2
31900 uppförandekoderna 1
31901 uppföranderegler 2
31902 uppförandereglerna 1
31903 uppförandet 3
31904 uppförde 2
31905 uppförs 1
31906 uppförstorad 1
31907 uppfört 1
31908 uppgavs 1
31909 uppger 1
31910 uppges 1
31911 uppgick 5
31912 uppgift 98
31913 uppgiften 9
31914 uppgifter 130
31915 uppgifterna 27
31916 uppgifternas 1
31917 uppgiftsfördelning 1
31918 uppgiftslämnare 1
31919 uppgiftsmängd 1
31920 uppgivande 1
31921 uppgradera 1
31922 uppgå 3
31923 uppgående 1
31924 uppgång 3
31925 uppgången 1
31926 uppgår 14
31927 uppgörelse 3
31928 uppgörelsen 2
31929 uppgörelser 2
31930 uppgörelserna 2
31931 upphandling 2
31932 upphetsad 1
31933 upphetsade 1
31934 upphetsande 1
31935 upphetsat 1
31936 upphetsning 1
31937 upphettat 1
31938 upphov 33
31939 upphovet 1
31940 upphovskällan 1
31941 upphovsman 4
31942 upphovsmannen 2
31943 upphovsmän 2
31944 upphovsmännen 4
31945 upphovsmännens 1
31946 upphovsrätt 11
31947 upphovsrätten 4
31948 upphovsrättsavgift 1
31949 upphovsrättsliga 1
31950 upphovsrättsligt 1
31951 upphovsrättsreglering 1
31952 upphängd 1
31953 upphängda 1
31954 upphäva 8
31955 upphävande 2
31956 upphävandet 3
31957 upphävas 5
31958 upphävdes 1
31959 upphävs 2
31960 upphöja 1
31961 upphöjda 2
31962 upphöjs 1
31963 upphör 7
31964 upphöra 14
31965 upphörandet 1
31966 upphörde 5
31967 upphört 7
31968 uppifrån 2
31969 uppkallad 1
31970 uppklädd 1
31971 uppkomma 2
31972 uppkommer 8
31973 uppkommit 5
31974 upplagan 1
31975 uppleva 14
31976 upplevde 5
31977 upplevelse 4
31978 upplevelser 1
31979 upplevelses 1
31980 upplever 14
31981 upplevs 2
31982 upplevt 6
31983 upplyftande 1
31984 upplysa 7
31985 upplyses 1
31986 upplysning 6
31987 upplysningar 5
31988 upplyst 7
31989 upplysta 1
31990 upplyste 2
31991 upplysts 1
31992 upplåsta 1
31993 upplösa 1
31994 upplöses 1
31995 upplösning 6
31996 upplösta 1
31997 upplöstes 2
31998 uppmana 28
31999 uppmanade 5
32000 uppmanades 1
32001 uppmanar 69
32002 uppmanas 12
32003 uppmanat 3
32004 uppmaning 11
32005 uppmaningar 3
32006 uppmaningen 2
32007 uppmaningsskrivelse 1
32008 uppmjukning 3
32009 uppmjukningen 2
32010 uppmuntra 37
32011 uppmuntrad 1
32012 uppmuntran 5
32013 uppmuntrande 9
32014 uppmuntrar 18
32015 uppmuntras 12
32016 uppmuntrat 2
32017 uppmuntrats 1
32018 uppmärksam 5
32019 uppmärksamhet 76
32020 uppmärksamheten 16
32021 uppmärksamma 23
32022 uppmärksammade 2
32023 uppmärksammar 4
32024 uppmärksammare 1
32025 uppmärksammas 7
32026 uppmärksammat 2
32027 uppmärksammats 1
32028 uppmärksamt 11
32029 uppmätta 1
32030 uppmättes 1
32031 uppnå 139
32032 uppnåbara 1
32033 uppnådda 6
32034 uppnådde 3
32035 uppnåddes 2
32036 uppnåeligt 1
32037 uppnår 21
32038 uppnås 36
32039 uppnått 20
32040 uppnåtts 17
32041 uppochner 1
32042 uppochnervända 1
32043 uppoffrande 1
32044 uppoffrat 1
32045 uppoffring 1
32046 uppoffringar 2
32047 upprensningar 1
32048 upprensningen 1
32049 upprepa 38
32050 upprepade 27
32051 upprepades 1
32052 upprepandets 1
32053 upprepar 41
32054 upprepas 15
32055 upprepat 4
32056 upprepats 3
32057 upprepning 2
32058 uppriktig 1
32059 uppriktiga 2
32060 uppriktighet 1
32061 uppriktigt 15
32062 upprivande 1
32063 upprop 2
32064 uppror 1
32065 upproriska 1
32066 upprusta 1
32067 uppryckning 1
32068 uppräknade 1
32069 uppräkning 2
32070 upprätta 29
32071 upprättade 2
32072 upprättades 1
32073 upprättande 4
32074 upprättandet 10
32075 upprättar 14
32076 upprättas 6
32077 upprättat 9
32078 upprättats 3
32079 upprättelse 1
32080 upprätthålla 20
32081 upprätthållande 1
32082 upprätthållandet 4
32083 upprätthållas 2
32084 upprätthåller 3
32085 upprätthållit 1
32086 upprätthålls 3
32087 uppröjningsarbetet 1
32088 uppröra 1
32089 upprörande 5
32090 uppröras 1
32091 upprörd 1
32092 upprörda 2
32093 upprördhet 1
32094 uppsamling 3
32095 uppsamlingen 1
32096 uppsamlingscentrum 1
32097 uppsamlingsplatser 2
32098 uppsamlingsplatserna 1
32099 uppsatt 4
32100 uppsatta 4
32101 uppseendeväckande 3
32102 uppsjö 1
32103 uppskakade 1
32104 uppskatta 7
32105 uppskattad 1
32106 uppskattade 4
32107 uppskattande 2
32108 uppskattar 22
32109 uppskattas 3
32110 uppskattat 1
32111 uppskattning 16
32112 uppskattningar 2
32113 uppskattningsvis 1
32114 uppskjuta 2
32115 uppskjutande 3
32116 uppskjutas 2
32117 uppskjuten 1
32118 uppskjuter 1
32119 uppskov 1
32120 uppskovet 1
32121 uppskruvade 3
32122 uppslagen 1
32123 uppslitsade 1
32124 uppsluppna 1
32125 uppsluppnaste 1
32126 uppslutning 1
32127 uppspaltning 1
32128 uppsplittring 1
32129 uppspärrade 1
32130 uppspårandet 1
32131 uppspårningsfasen 1
32132 uppstaplade 1
32133 uppstod 8
32134 uppsträckta 1
32135 uppströms 5
32136 uppställa 2
32137 uppställandet 1
32138 uppställas 1
32139 uppställda 5
32140 uppställer 1
32141 uppställning 1
32142 uppställningsspår 1
32143 uppstå 17
32144 uppståndelse 1
32145 uppståndelsen 1
32146 uppstår 47
32147 uppstått 19
32148 uppsving 5
32149 uppsyn 1
32150 uppsägning 1
32151 uppsägningar 11
32152 uppsägningsbesked 1
32153 uppsägningsbeskedet 1
32154 uppsättning 4
32155 upptagen 5
32156 upptaget 4
32157 upptagetton 1
32158 upptagit 1
32159 upptagits 1
32160 upptagna 2
32161 upptagningsområde 1
32162 upptar 3
32163 upptas 3
32164 upptrappningen 1
32165 uppträda 2
32166 uppträdande 9
32167 uppträdde 1
32168 uppträder 8
32169 uppträtt 1
32170 upptäcka 7
32171 upptäcker 6
32172 upptäcks 3
32173 upptäckt 6
32174 upptäckte 17
32175 upptäckten 3
32176 upptäcktes 3
32177 upptäckts 5
32178 upptäcktsfärdernas 1
32179 uppvaknad 1
32180 uppviglande 1
32181 uppvisa 5
32182 uppvisade 1
32183 uppvisar 11
32184 uppvisas 1
32185 uppvisat 4
32186 uppväga 3
32187 uppväger 1
32188 uppvända 1
32189 uppvärdera 1
32190 uppvärderar 2
32191 uppvärdering 2
32192 uppäten 1
32193 uppåt 8
32194 ur 143
32195 uran 8
32196 uranium 2
32197 uranvapen 4
32198 urartad 1
32199 urartade 1
32200 urartande 1
32201 urartar 1
32202 urban 3
32203 urbana 4
32204 urbanisering 1
32205 urbaniseringen 2
32206 urgamla 1
32207 urgammal 1
32208 urholka 3
32209 urholkar 1
32210 urholkas 4
32211 urholkat 1
32212 urholkningen 1
32213 urminnes 1
32214 urringning 1
32215 ursinnig 1
32216 urskilja 5
32217 urskiljas 1
32218 urskiljer 3
32219 urskillningslöst 1
32220 urskogar 1
32221 urskuldande 1
32222 ursprung 25
32223 ursprunget 6
32224 ursprungliga 47
32225 ursprungligen 9
32226 ursprungsbefolkning 1
32227 ursprungsbefolkningar 4
32228 ursprungsbestämmelser 1
32229 ursprungsfrågor 1
32230 ursprungsintyg 1
32231 ursprungskick 1
32232 ursprungsland 2
32233 ursprungslandet 1
32234 ursprungsländer 1
32235 ursprungsländerna 3
32236 ursprungsmärkning 1
32237 ursprungsregionerna 1
32238 ursprungsregler 2
32239 ursprungsreglerna 1
32240 ursprungsversionen 1
32241 urspårning 1
32242 ursäkt 20
32243 ursäkta 9
32244 ursäktade 1
32245 ursäktande 2
32246 ursäkten 2
32247 ursäkter 4
32248 urtider 1
32249 urval 5
32250 urvalet 5
32251 urvalsfråga 2
32252 urvalsfrågan 1
32253 urvalskommittéerna 1
32254 urvalskriterier 2
32255 urvalskriterierna 2
32256 urvattna 2
32257 urvattnade 1
32258 urvattnar 2
32259 urvattnas 3
32260 urvattnat 1
32261 urvattning 3
32262 uråldriga 1
32263 uråldrigare 1
32264 ut 491
32265 ut-och-invändningsteknik 1
32266 utan 935
32267 utanför 104
32268 utanförskap 3
32269 utanpå 1
32270 utantill 1
32271 utarbeta 42
32272 utarbetade 6
32273 utarbetades 3
32274 utarbetande 1
32275 utarbetandet 19
32276 utarbetar 9
32277 utarbetas 9
32278 utarbetat 9
32279 utarbetats 6
32280 utarmade 5
32281 utarmar 1
32282 utarmas 1
32283 utarmat 6
32284 utarmningen 1
32285 utbasunerade 1
32286 utbetalade 3
32287 utbetalades 1
32288 utbetalas 1
32289 utbetalning 3
32290 utbetalningar 1
32291 utbetalningarna 1
32292 utbetalningen 2
32293 utbilda 4
32294 utbildade 4
32295 utbildar 2
32296 utbildas 4
32297 utbildats 1
32298 utbildning 63
32299 utbildningar 2
32300 utbildningen 9
32301 utbildningens 1
32302 utbildnings- 5
32303 utbildningscentra 1
32304 utbildningscentren 1
32305 utbildningsinsatser 1
32306 utbildningsinstitutioner 2
32307 utbildningskostnader 2
32308 utbildningsministern 1
32309 utbildningsmoment 1
32310 utbildningsmöjligheter 1
32311 utbildningsnivå 3
32312 utbildningsnivån 1
32313 utbildningsoffensiv 1
32314 utbildningsområdet 1
32315 utbildningspolitiken 2
32316 utbildningspolitisk 2
32317 utbildningspraktik 1
32318 utbildningsprogram 2
32319 utbildningsprojekt 1
32320 utbildningssamhälle 1
32321 utbildningsstrukturer 1
32322 utbildningssystem 1
32323 utbildningssystemens 1
32324 utbildningssystemet 1
32325 utbildningsåtgärder 1
32326 utblottade 1
32327 utbrast 1
32328 utbredd 3
32329 utbredda 1
32330 utbredning 6
32331 utbredningen 1
32332 utbrister 1
32333 utbrott 3
32334 utbrottet 1
32335 utbrutit 1
32336 utbrytarstyrkor 1
32337 utbud 6
32338 utbudet 2
32339 utbudsinriktad 1
32340 utbyggd 1
32341 utbyggnad 4
32342 utbyggnaden 2
32343 utbyggt 1
32344 utbyta 4
32345 utbyte 30
32346 utbyten 1
32347 utbyter 2
32348 utbytesprincipen 1
32349 utbytesprojekt 2
32350 utbytet 6
32351 utbytte 2
32352 utbärningar 1
32353 utdela 1
32354 utdelad 1
32355 utdelar 1
32356 utdelas 2
32357 utdelning 3
32358 utdelningen 2
32359 utdrag 1
32360 utdragen 2
32361 utdragna 2
32362 utdömda 1
32363 utdömer 2
32364 ute 35
32365 uteblivit 1
32366 utedasset 1
32367 utefter 1
32368 utelämna 1
32369 utelämnade 1
32370 utelämnas 4
32371 utesluta 6
32372 uteslutande 15
32373 uteslutas 2
32374 utesluten 1
32375 utesluter 7
32376 uteslutet 2
32377 uteslutits 1
32378 uteslutna 1
32379 uteslutning 6
32380 utesluts 1
32381 uteslöt 2
32382 utestänga 1
32383 utestängas 4
32384 utestängda 1
32385 utestängning 2
32386 utestängs 1
32387 utestängt 1
32388 utestängts 1
32389 utfall 1
32390 utfallet 1
32391 utfarten 1
32392 utfasning 3
32393 utfasningen 4
32394 utfiskning 1
32395 utflaggningsländer 1
32396 utflykter 2
32397 utflyttade 1
32398 utflyttningen 1
32399 utflyttningsbidrag 1
32400 utfodrat 1
32401 utforma 24
32402 utformad 2
32403 utformade 9
32404 utformades 1
32405 utformandet 3
32406 utformar 6
32407 utformas 13
32408 utformat 4
32409 utformats 1
32410 utformning 21
32411 utformningar 1
32412 utformningen 21
32413 utformningsmässiga 1
32414 utforska 2
32415 utforskas 1
32416 utfrågning 9
32417 utfrågningar 1
32418 utfrågningarna 1
32419 utfrågningen 4
32420 utfärda 8
32421 utfärdades 1
32422 utfärdande 4
32423 utfärdandet 2
32424 utfärdar 1
32425 utfärdas 1
32426 utfärdat 3
32427 utfärdats 1
32428 utfästelser 2
32429 utför 13
32430 utföra 28
32431 utförande 2
32432 utföras 2
32433 utförd 1
32434 utförda 2
32435 utförde 2
32436 utfördes 2
32437 utförlig 2
32438 utförliga 2
32439 utförligare 1
32440 utförligen 1
32441 utförligt 2
32442 utförs 8
32443 utfört 13
32444 utförts 6
32445 utgallring 4
32446 utgallringen 1
32447 utgavs 1
32448 utgick 3
32449 utgifter 27
32450 utgifterna 11
32451 utgifts 1
32452 utgiftsmål 1
32453 utgiftsområde 11
32454 utgiftsområden 1
32455 utgiftsområdet 1
32456 utgiftspolitik 1
32457 utgiftsprioriteringar 1
32458 utgiftsprogram 1
32459 utgiftssektorer 1
32460 utgiftstak 1
32461 utgivare 1
32462 utgivit 1
32463 utgivna 2
32464 utgjorde 10
32465 utgjordes 1
32466 utgjort 3
32467 utgrävningen 1
32468 utgå 11
32469 utgång 4
32470 utgången 9
32471 utgångsförslag 1
32472 utgångsläge 1
32473 utgångspunkt 22
32474 utgångspunkten 5
32475 utgångspunkter 4
32476 utgår 25
32477 utgått 4
32478 utgåva 1
32479 utgåvor 1
32480 utgör 135
32481 utgöra 34
32482 utgörs 8
32483 utgör­ 1
32484 uthuset 1
32485 uthyrning 5
32486 uthärda 1
32487 uthärdliga 1
32488 uthållighet 2
32489 utifrån 48
32490 utjämna 4
32491 utjämningen 1
32492 utjämningsfond 1
32493 utkanten 4
32494 utkast 13
32495 utkasten 1
32496 utkastet 10
32497 utkik 1
32498 utkom 1
32499 utkomst 3
32500 utkonkurrerade 1
32501 utkräva 1
32502 utkrävandet 1
32503 utkräver 2
32504 utkämpa 2
32505 utkämpar 1
32506 utlandet 4
32507 utlandsplacerade 2
32508 utlandsplacering 1
32509 utloppet 1
32510 utlovade 7
32511 utlovar 1
32512 utlovat 3
32513 utlovats 1
32514 utlyst 2
32515 utlägg 1
32516 utläggningar 1
32517 utlämna 1
32518 utlämnad 1
32519 utlämnats 1
32520 utlämning 1
32521 utländsk 2
32522 utländska 10
32523 utlänningslagarna 1
32524 utlänningslagen 2
32525 utläsa 1
32526 utlåning 2
32527 utlåtande 1
32528 utlåtanden 1
32529 utlåtandet 1
32530 utlösa 1
32531 utlösande 1
32532 utlöst 1
32533 utlöste 1
32534 utlöstes 1
32535 utmana 3
32536 utmanande 3
32537 utmanas 1
32538 utmaning 31
32539 utmaningar 36
32540 utmaningarna 7
32541 utmaningen 15
32542 utmattning 1
32543 utmed 4
32544 utmynnar 1
32545 utmynnat 1
32546 utmärkande 1
32547 utmärker 3
32548 utmärks 2
32549 utmärkt 46
32550 utmärkta 38
32551 utnyttja 56
32552 utnyttjade 2
32553 utnyttjades 3
32554 utnyttjande 14
32555 utnyttjandet 7
32556 utnyttjar 11
32557 utnyttjas 19
32558 utnyttjat 5
32559 utnyttjats 1
32560 utnämna 3
32561 utnämnandet 1
32562 utnämndes 1
32563 utnämner 1
32564 utnämning 1
32565 utnämningen 1
32566 utnämnt 1
32567 utnämnts 2
32568 utom 12
32569 utomeuropeiska 6
32570 utomeuropeiskt 1
32571 utomhus 1
32572 utomlands 2
32573 utomordentlig 1
32574 utomordentliga 3
32575 utomordentligt 16
32576 utomstående 5
32577 utopier 1
32578 utopiskt 1
32579 utpeka 1
32580 utpekar 1
32581 utpekas 1
32582 utplacerad 1
32583 utplacerade 2
32584 utplacerades 1
32585 utplacering 2
32586 utplåna 4
32587 utplånade 1
32588 utplånande 1
32589 utplånar 1
32590 utplånat 1
32591 utplåning 3
32592 utpressning 3
32593 utpräglad 1
32594 utpräglade 1
32595 utrangeras 1
32596 utreda 3
32597 utredande 2
32598 utredd 1
32599 utredning 4
32600 utredningar 5
32601 utredningarna 1
32602 utredningsarbetet 1
32603 utredningsbyråer 1
32604 utredningshäktning 1
32605 utredningstekniska 1
32606 utredningsverksamhet 1
32607 utreds 1
32608 utrikes 3
32609 utrikes- 20
32610 utrikesdepartementet 2
32611 utrikesenhet 1
32612 utrikesfrågor 13
32613 utrikesförbindelser 2
32614 utrikeshandel 5
32615 utrikeshandelspolitikerna 1
32616 utrikeskorrespondenter 1
32617 utrikesminister 3
32618 utrikesministeriernas 1
32619 utrikesministern 7
32620 utrikesministrarna 2
32621 utrikesnivå 1
32622 utrikespolitik 12
32623 utrikespolitiken 15
32624 utrikespolitisk 1
32625 utrikespolitiska 4
32626 utropa 1
32627 utropar 1
32628 utropas 2
32629 utrota 16
32630 utrotad 1
32631 utrotas 2
32632 utrotning 2
32633 utrotningar 1
32634 utrotningen 2
32635 utrotningshotade 1
32636 utrotningsstrategier 1
32637 utrotningsåtgärder 1
32638 utrullad 1
32639 utrustad 1
32640 utrustade 1
32641 utrustar 2
32642 utrustas 2
32643 utrustning 8
32644 utrustningar 1
32645 utrustningen 2
32646 utrymme 23
32647 utrymmet 1
32648 uträtta 6
32649 uträttar 1
32650 uträttat 2
32651 utröna 3
32652 utsatt 5
32653 utsatta 10
32654 utsattes 1
32655 utsatthet 1
32656 utsatts 3
32657 utse 4
32658 utsedd 1
32659 utsedda 2
32660 utseende 9
32661 utser 2
32662 utses 3
32663 utsett 2
32664 utsetts 1
32665 utsikt 3
32666 utsikten 3
32667 utsikter 3
32668 utsikterna 5
32669 utsirade 1
32670 utskott 59
32671 utskotten 7
32672 utskottet 290
32673 utskottets 16
32674 utskotts 3
32675 utskottsbehandlingen 5
32676 utskottsdebatten 1
32677 utskottsförhandlingen 1
32678 utskottsrummen 1
32679 utskottssammanträdet 1
32680 utskottssekretariatet 1
32681 utslag 3
32682 utslagen 1
32683 utslagna 4
32684 utslagning 20
32685 utslagningen 6
32686 utslagningens 1
32687 utslagningsmekanismer 1
32688 utslagningspolitik 1
32689 utslungade 1
32690 utsläpp 15
32691 utsläppen 11
32692 utsläppet 5
32693 utsläppsnivåer 1
32694 utsläppsrätter 1
32695 utslätning 1
32696 utspelad 1
32697 utspelade 2
32698 utspridd 1
32699 utspridda 2
32700 utspridning 1
32701 utspärrade 1
32702 utstationera 1
32703 utstationerad 1
32704 utstationerade 1
32705 utstationering 7
32706 utstationeringssituationen 1
32707 utsträcka 1
32708 utsträckas 2
32709 utsträckning 69
32710 utsträckningen 1
32711 utsträcks 1
32712 utsträckt 1
32713 utsträckta 1
32714 utstrålade 1
32715 utstrålar 1
32716 utströdda 1
32717 utstuderad 1
32718 utställandet 1
32719 utställda 1
32720 utställningar 4
32721 utställningsföremål 1
32722 utställt 1
32723 utstå 5
32724 utstående 2
32725 utstår 1
32726 utstått 2
32727 utstötta 3
32728 utsugare 2
32729 utsugning 1
32730 utsvulten 1
32731 utsäde 4
32732 utsända 1
32733 utsätta 6
32734 utsättas 5
32735 utsätter 1
32736 utsättningsdirektivet 1
32737 utsätts 11
32738 utsågs 3
32739 utsålda 1
32740 utsökta 1
32741 uttag 1
32742 uttagningsprov 1
32743 uttala 38
32744 uttalad 3
32745 uttalade 17
32746 uttalades 3
32747 uttalande 89
32748 uttalanden 47
32749 uttalandena 4
32750 uttalandet 10
32751 uttalar 17
32752 uttalas 4
32753 uttalat 17
32754 uttaxeraren 1
32755 uttjänta 25
32756 uttolkare 1
32757 uttolkarna 1
32758 uttorkning 2
32759 uttrar 1
32760 uttryck 67
32761 uttrycka 48
32762 uttryckas 1
32763 uttrycker 13
32764 uttrycket 9
32765 uttrycklig 2
32766 uttryckliga 3
32767 uttryckligen 20
32768 uttryckligt 1
32769 uttrycks 13
32770 uttrycksfull 1
32771 uttryckslös 1
32772 uttryckt 16
32773 uttryckta 2
32774 uttryckte 19
32775 uttrycktes 3
32776 uttryckts 4
32777 utträda 1
32778 utträde 1
32779 uttänkt 1
32780 uttänkta 1
32781 uttömd 1
32782 uttömda 1
32783 uttömmande 6
32784 uttömt 1
32785 utvald 1
32786 utvalda 2
32787 utvandring 2
32788 utveckla 77
32789 utvecklad 4
32790 utvecklade 32
32791 utvecklades 2
32792 utvecklande 2
32793 utvecklandet 3
32794 utvecklar 8
32795 utvecklare 3
32796 utvecklaren 3
32797 utvecklas 59
32798 utvecklat 9
32799 utvecklats 12
32800 utveckling 284
32801 utvecklingar 1
32802 utvecklingen 168
32803 utvecklingens 2
32804 utvecklings- 9
32805 utvecklingsaktörer 1
32806 utvecklingsarbete 1
32807 utvecklingsaspekterna 1
32808 utvecklingsbistånd 7
32809 utvecklingsbiståndet 1
32810 utvecklingsbiståndsprogram 1
32811 utvecklingsbudget 1
32812 utvecklingscentrum 1
32813 utvecklingscentrumet 1
32814 utvecklingsfas 2
32815 utvecklingsfond 1
32816 utvecklingsfonden 15
32817 utvecklingsfondens 1
32818 utvecklingsfonder 1
32819 utvecklingsfrämjande 1
32820 utvecklingsfråga 2
32821 utvecklingsfrågan 1
32822 utvecklingsfrågor 3
32823 utvecklingsfunktioner 1
32824 utvecklingsfunktionerna 1
32825 utvecklingsförmåga 1
32826 utvecklingshjälp 1
32827 utvecklingshjälpen 1
32828 utvecklingsinitiativ 1
32829 utvecklingsinsatser 1
32830 utvecklingsinstrument 1
32831 utvecklingskonferens 1
32832 utvecklingsland 1
32833 utvecklingsländer 15
32834 utvecklingsländerna 42
32835 utvecklingsländernas 7
32836 utvecklingsmetod 1
32837 utvecklingsminister 1
32838 utvecklingsmodell 2
32839 utvecklingsmässigt 1
32840 utvecklingsmål 1
32841 utvecklingsmålen 3
32842 utvecklingsmöjligheter 1
32843 utvecklingsmöjligheterna 1
32844 utvecklingsmönster 1
32845 utvecklingsnationerna 2
32846 utvecklingsnivå 1
32847 utvecklingsnivåer 2
32848 utvecklingsområde 1
32849 utvecklingsområden 1
32850 utvecklingsområdet 3
32851 utvecklingspartner 2
32852 utvecklingspartnerskap 4
32853 utvecklingspartnerskapen 1
32854 utvecklingspartnerskapens 1
32855 utvecklingsperspektivet 1
32856 utvecklingsplan 1
32857 utvecklingsplanerna 1
32858 utvecklingspolicy 1
32859 utvecklingspolitik 14
32860 utvecklingspolitiken 36
32861 utvecklingspotential 1
32862 utvecklingsprioriteringar 1
32863 utvecklingsprioriteringarna 1
32864 utvecklingsprocess 2
32865 utvecklingsprocessen 1
32866 utvecklingsprogram 4
32867 utvecklingsprogrammen 6
32868 utvecklingsprojekt 2
32869 utvecklingsprojekten 1
32870 utvecklingsprojekts 1
32871 utvecklingsredskapet 1
32872 utvecklingssamarbete 9
32873 utvecklingssamarbetesaspekten 1
32874 utvecklingssamarbetet 5
32875 utvecklingssamhället 1
32876 utvecklingsstadiet 2
32877 utvecklingssteg 1
32878 utvecklingsstrategi 1
32879 utvecklingsstrategier 3
32880 utvecklingsstrategierna 1
32881 utvecklingsstöd 6
32882 utvecklingsstödet 1
32883 utvecklingstakten 1
32884 utvecklingstjänstemän 1
32885 utvecklingstjänsterna 1
32886 utvecklingsväg 1
32887 utvecklingsändamål 1
32888 utverka 5
32889 utvidga 28
32890 utvidgad 5
32891 utvidgade 3
32892 utvidgades 1
32893 utvidgande 1
32894 utvidgar 8
32895 utvidgas 18
32896 utvidgat 3
32897 utvidgning 49
32898 utvidgningar 2
32899 utvidgningarna 1
32900 utvidgningen 99
32901 utvidgningens 4
32902 utvidgningsfrågan 1
32903 utvidgningsplanerna 1
32904 utvidgningsprocess 1
32905 utvidgningsprocessen 6
32906 utvidgningsprojektet 2
32907 utvidgningsrunda 1
32908 utvidgningsärendet 1
32909 utvinningsnivåer 1
32910 utvinns 1
32911 utvisa 3
32912 utvisade 1
32913 utvisar 1
32914 utvisning 3
32915 utväg 4
32916 utvärdera 12
32917 utvärderar 2
32918 utvärderas 6
32919 utvärderat 1
32920 utvärdering 30
32921 utvärderingar 6
32922 utvärderingarna 1
32923 utvärderingen 15
32924 utvärderingskommittéerna 1
32925 utvärderingspanelerna 1
32926 utväxlade 2
32927 utväxlandet 1
32928 utväxlat 1
32929 utväxling 2
32930 utåt 5
32931 utöka 13
32932 utökad 2
32933 utökade 1
32934 utökades 2
32935 utökande 1
32936 utökar 2
32937 utökas 4
32938 utökat 3
32939 utökning 2
32940 utöva 18
32941 utövade 1
32942 utövades 1
32943 utövande 8
32944 utövandet 2
32945 utövar 9
32946 utövas 9
32947 utövat 1
32948 utöver 24
32949 v 1
32950 va 3
32951 vaccin 10
32952 vaccination 2
32953 vaccinationsprogram 1
32954 vacciner 1
32955 vaccinera 1
32956 vaccinering 5
32957 vaccinet 1
32958 vacker 8
32959 vackert 2
32960 vackla 1
32961 vackra 23
32962 vackraste 2
32963 vad 735
32964 vag 1
32965 vaga 11
32966 vagabond 1
32967 vaggan 1
32968 vagnar 1
32969 vagnen 3
32970 vagt 3
32971 vajande 1
32972 vaka 2
32973 vakande 1
32974 vakar 2
32975 vaken 1
32976 vaket 1
32977 vakna 2
32978 vaknade 7
32979 vaknar 2
32980 vaksam 6
32981 vaksamhet 4
32982 vaksamma 10
32983 vaksammare 1
32984 vaksamt 2
32985 vakt 3
32986 vakter 1
32987 vaktmästarna 1
32988 vakuum 3
32989 vakuumtankar 1
32990 val 46
32991 valbarhet 1
32992 valbart 1
32993 vald 10
32994 valda 19
32995 valdagen 1
32996 valde 6
32997 valdeltagandet 7
32998 valdes 4
32999 valdistrikt 2
33000 valen 10
33001 valet 17
33002 valfläsk 1
33003 valframgång 1
33004 valframgångar 2
33005 valfrihet 1
33006 valfriheten 2
33007 valfråga 1
33008 valfusket 1
33009 valförfaranden 1
33010 valkampanj 3
33011 valkampanjen 2
33012 valkampanjerna 1
33013 valkrets 6
33014 valkretsar 1
33015 valkretsen 1
33016 vallfärd 1
33017 vallfärdsstav 1
33018 vallistorna 2
33019 vallokalerna 1
33020 valmässiga 1
33021 valmöjligheter 2
33022 valnötsträden 1
33023 valobservation 1
33024 valobservatörer 1
33025 valområden 1
33026 valperioden 1
33027 valresultaten 1
33028 valresultatet 2
33029 valrörelse 1
33030 valrörelsen 1
33031 valsedlar 1
33032 valseger 1
33033 valt 19
33034 valtaktiska 1
33035 valtider 2
33036 valts 9
33037 valuation 1
33038 valuta 18
33039 valutafonden 4
33040 valutafondens 1
33041 valutafrågor 27
33042 valutaförfalskare 1
33043 valutaförfalskning 3
33044 valutaförfalskningar 1
33045 valutaförfalskningen 1
33046 valutaförfalskningsbrott 1
33047 valutan 21
33048 valutans 4
33049 valutapolitikens 1
33050 valutarisker 1
33051 valutaspekulationen 2
33052 valutaunionen 3
33053 valutaunionens 1
33054 valutor 5
33055 valutorna 3
33056 valv 2
33057 valven 1
33058 valörer 1
33059 valövervakningen 1
33060 vampyr 1
33061 van 38
33062 vana 4
33063 vandra 5
33064 vandrade 6
33065 vandrande 1
33066 vandrare 1
33067 vandringar 1
33068 vanhedra 1
33069 vanhedrande 2
33070 vanlig 11
33071 vanliga 21
33072 vanligare 5
33073 vanligaste 3
33074 vanligen 2
33075 vanligt 14
33076 vanligtvis 5
33077 vann 3
33078 vanor 3
33079 vansinne 3
33080 vansinnig 1
33081 vansinnigheter 1
33082 vansklig 1
33083 vanskliga 2
33084 vapen 22
33085 vapendragaren 1
33086 vapenhandeln 2
33087 vapenhandlare 1
33088 vapenindustrin 1
33089 vapenolja 1
33090 vapenrocken 1
33091 vapenvila 2
33092 vapenvilan 1
33093 vapnen 3
33094 var 1182
33095 vara 1159
33096 varade 2
33097 varaktig 10
33098 varaktiga 4
33099 varaktigt 4
33100 varan 3
33101 varandra 82
33102 varandras 3
33103 varann 1
33104 varannan 1
33105 varans 1
33106 varat 3
33107 varav 10
33108 varböld 2
33109 vardag 2
33110 vardagar 1
33111 vardagen 3
33112 vardagliga 5
33113 vardagligt 3
33114 vardags 1
33115 vardagsfraser 1
33116 vardagskriminaliteten 1
33117 vardagslag 1
33118 vardagsmat 1
33119 vardagspolitiken 1
33120 vardagsrum 1
33121 vardagsrummet 8
33122 vardagsrutin 1
33123 vardande 1
33124 vardera 1
33125 vare 100
33126 varefter 6
33127 varelse 2
33128 varelsen 1
33129 varelser 3
33130 varelserna 1
33131 varenda 16
33132 varför 114
33133 vargar 1
33134 vargarna 2
33135 varhelst 3
33136 vari 2
33137 variabel 2
33138 variabler 2
33139 variant 1
33140 varianter 1
33141 varierade 1
33142 varierande 4
33143 varierar 5
33144 varierat 1
33145 varifrån 5
33146 varigenom 2
33147 varit 304
33148 varje 276
33149 varken 47
33150 varm 3
33151 varma 9
33152 varmaste 1
33153 varmblodiga 1
33154 varmed 1
33155 varmt 27
33156 varmvattenberedaren 1
33157 varna 7
33158 varnade 2
33159 varnades 1
33160 varnagel 1
33161 varnande 1
33162 varnar 4
33163 varnat 2
33164 varning 14
33165 varningar 1
33166 varningarna 1
33167 varningen 1
33168 varningens 1
33169 varningssignal 1
33170 varningssystemet 1
33171 varor 20
33172 varorna 3
33173 varors 2
33174 varpbomtrålare 1
33175 varpå 4
33176 vars 83
33177 varsamma 1
33178 varse 1
33179 varsel 3
33180 varslar 1
33181 varstans 1
33182 varsågod 1
33183 vart 25
33184 vartannat 4
33185 vartenda 2
33186 varv 2
33187 varvid 12
33188 varvsindustrin 2
33189 varvsstöd 2
33190 vaska 1
33191 vassa 1
33192 vatten 127
33193 vatten- 1
33194 vattenanvändarna 4
33195 vattenanvändning 4
33196 vattenanvändningen 1
33197 vattenavgifter 3
33198 vattenbrist 6
33199 vattenbruk 5
33200 vattenbruket 2
33201 vattenbrukets 1
33202 vattenbruksanläggningar 1
33203 vattenbruksindustrin 2
33204 vattenbruksnäringen 1
33205 vattenbrukssektorn 4
33206 vattenbrukssystem 1
33207 vattenbrukssystemen 1
33208 vattenbyggnadsarbeten 1
33209 vattendammar 1
33210 vattendelare 2
33211 vattendirektiv 1
33212 vattendirektivet 2
33213 vattendistributionen 1
33214 vattendrag 5
33215 vattendragen 2
33216 vattendunkar 1
33217 vattenekosystem 1
33218 vattenextraktion 1
33219 vattenflöde 1
33220 vattenfrågan 1
33221 vattenfylld 1
33222 vattenfördelningen 1
33223 vattenföroreningar 1
33224 vattenförråden 1
33225 vattenförsämring 2
33226 vattenförsörjning 1
33227 vattenförsörjningen 1
33228 vattenförvaltning 1
33229 vattenförvaltningen 1
33230 vattengränser 1
33231 vattenhushållning 2
33232 vattenindikatorerna 1
33233 vattenkatastrof 1
33234 vattenkostnaden 1
33235 vattenkostnaderna 1
33236 vattenkraftsprojekt 1
33237 vattenkrig 1
33238 vattenkvalitet 6
33239 vattenkvaliteten 5
33240 vattenkvalitetområden 1
33241 vattenkällorna 1
33242 vattenlagstiftning 1
33243 vattenlagstiftningen 1
33244 vattenleverantörerna 1
33245 vattenmiljö 1
33246 vattenmiljön 6
33247 vattenmyndigheter 1
33248 vattenmyndigheterna 1
33249 vattenmängden 1
33250 vattenmätare 1
33251 vattennyttjande 1
33252 vattennät 1
33253 vattenområde 1
33254 vattenområden 3
33255 vattenområdet 2
33256 vattenpolitik 8
33257 vattenpolitiken 11
33258 vattenpolitikens 6
33259 vattenpriser 1
33260 vattenprispolitiken 1
33261 vattenproblematiken 1
33262 vattenproblemen 1
33263 vattenramdirektivet 1
33264 vattenramdirektivets 1
33265 vattenrening 1
33266 vattenreningsanläggningar 1
33267 vattenreningsutrustning 1
33268 vattenreserver 2
33269 vattenreserverna 2
33270 vattenreservernas 1
33271 vattenresurser 6
33272 vattenresurserna 12
33273 vattensaneringen 1
33274 vattensituation 1
33275 vattenskydd 1
33276 vattenskyddet 2
33277 vattenskyddslagstiftning 1
33278 vattenslöseri 1
33279 vattensystem 2
33280 vattensystemen 1
33281 vattensystemet 2
33282 vattentermer 1
33283 vattenterritorium 1
33284 vattentillgångar 1
33285 vattentillgången 1
33286 vattenutnyttjande 6
33287 vattenväg 2
33288 vattenvägar 8
33289 vattenvården 1
33290 vattenöverflöd 1
33291 vattnade 1
33292 vattnas 1
33293 vattnen 1
33294 vattnet 62
33295 vattnets 3
33296 veck 1
33297 vecka 24
33298 veckan 42
33299 veckans 1
33300 veckas 1
33301 veckobesök 1
33302 veckor 35
33303 veckorna 17
33304 veckoslut 1
33305 veckosluten 1
33306 veckotidningar 1
33307 ved 3
33308 vederbörande 2
33309 vederbörandes 1
33310 vederbörlig 10
33311 vederbörliga 2
33312 vederbörligen 4
33313 vederbörligt 3
33314 vedergällningsaktion 1
33315 vederkvickande 1
33316 vederlägger 1
33317 vedermödor 1
33318 vedertagna 1
33319 vedervärdiga 1
33320 vek 3
33321 vekhet 3
33322 vekheten 1
33323 velat 21
33324 vem 59
33325 vems 2
33326 ventileras 1
33327 ventures 1
33328 veranda 1
33329 verandan 2
33330 verbala 1
33331 verifiable 1
33332 verifierbara 1
33333 verk 12
33334 verka 25
33335 verkade 23
33336 verkan 9
33337 verkar 112
33338 verkat 4
33339 verket 77
33340 verkets 2
33341 verklig 61
33342 verkliga 72
33343 verklige 1
33344 verkligen 342
33345 verklighet 29
33346 verkligheten 48
33347 verkligheterna 1
33348 verklighetsfrämmande 1
33349 verkligt 52
33350 verkningar 1
33351 verkningsfulla 1
33352 verkningsfullt 4
33353 verkningslösa 2
33354 verkningslöst 2
33355 verksam 2
33356 verksamhet 93
33357 verksamheten 25
33358 verksamheter 11
33359 verksamheterna 2
33360 verksamhets 1
33361 verksamhetsavbrottet 1
33362 verksamhetsbas 1
33363 verksamhetsbudgetering 1
33364 verksamhetsgrenar 2
33365 verksamhetsmiljön 1
33366 verksamhetsområde 5
33367 verksamhetsprogram 1
33368 verksamhetstiden 1
33369 verksamhetstillväxt 1
33370 verksamhetsutveckling 1
33371 verksamhetsutövare 2
33372 verksamhetsutövarna 1
33373 verksamhetsutövarnas 1
33374 verksamhetsår 1
33375 verksamma 9
33376 verksamt 2
33377 verkstad 1
33378 verkstadsindustrin 1
33379 verkställa 7
33380 verkställande 9
33381 verkställandet 6
33382 verkställare 1
33383 verkställas 4
33384 verkställdes 1
33385 verkställer 3
33386 verkställighet 3
33387 verkställigheten 5
33388 verkställighetssynpunkt 1
33389 verkställs 2
33390 verkställts 1
33391 verktyg 18
33392 verktygen 1
33393 verktygsfält 1
33394 verktygsfältet 1
33395 verktygsstålstillverkarna 1
33396 versa 1
33397 versaler 3
33398 version 10
33399 versionen 16
33400 versioner 2
33401 versionsnumret 1
33402 vertikal 2
33403 vertikala 4
33404 vet 357
33405 veta 88
33406 vetat 2
33407 vetenskap 18
33408 vetenskapen 9
33409 vetenskapens 2
33410 vetenskaplig 20
33411 vetenskapliga 53
33412 vetenskapligt 8
33413 vetenskapsmän 11
33414 vetenskapsmännen 8
33415 vetenskapsmännens 1
33416 veteran- 1
33417 veteranbilar 6
33418 veteranbilarna 1
33419 veterinärer 1
33420 veterinärfrågor 1
33421 veterinärpersonal 1
33422 veterligen 1
33423 veto 6
33424 vetorätt 3
33425 vetoröster 1
33426 vetskap 3
33427 vetskapen 3
33428 vette 1
33429 vetter 3
33430 vettet 1
33431 vettig 5
33432 vettiga 1
33433 vettigt 5
33434 vettlös 1
33435 vettvilling 1
33436 vevade 1
33437 vi 4650
33438 via 55
33439 vibrerande 1
33440 vice 33
33441 vicelehendakari 1
33442 vicepresident 1
33443 vickade 1
33444 vid 629
33445 vida 9
33446 vidare 103
33447 vidarebefordra 5
33448 vidarebefordrar 1
33449 vidarebefordras 2
33450 vidarebefordrats 1
33451 vidarebehandlas 1
33452 vidareutbildning 1
33453 vidareutveckla 2
33454 vidareutvecklas 1
33455 vidareutvecklat 1
33456 vidareutveckling 1
33457 vidareutvecklingen 1
33458 vidaste 2
33459 vidbrättade 1
33460 vidd 2
33461 vidden 5
33462 video 1
33463 videoförhör 1
33464 videokonferenser 4
33465 vidga 2
33466 vidgades 2
33467 vidgas 1
33468 vidgå 1
33469 vidhålla 1
33470 vidhåller 4
33471 vidhållit 1
33472 vidhålls 1
33473 vidhöll 1
33474 vidmakthålla 3
33475 vidmakthållas 1
33476 vidriga 1
33477 vidröras 1
33478 vidrörd 1
33479 vidrörde 1
33480 vidskeplighet 1
33481 vidsträckt 1
33482 vidsynta 1
33483 vidta 93
33484 vidtaga 1
33485 vidtagit 10
33486 vidtagits 6
33487 vidtagna 4
33488 vidtalat 1
33489 vidtar 17
33490 vidtas 36
33491 vidtog 1
33492 vidtogs 5
33493 viftade 1
33494 viftades 1
33495 viftar 1
33496 vigt 1
33497 vigvattnet 1
33498 vigör 1
33499 vika 2
33500 vikarierna 1
33501 viker 2
33502 vikt 47
33503 vikt- 3
33504 vikten 24
33505 vikter 1
33506 viktförlust 1
33507 viktgränsen 2
33508 viktig 222
33509 viktiga 196
33510 viktigare 30
33511 viktigast 4
33512 viktigaste 124
33513 viktigt 401
33514 viktklasser 1
33515 vila 6
33516 vilade 2
33517 vilande 1
33518 vilar 19
33519 vilat 1
33520 vild 4
33521 vilda 14
33522 vildar 1
33523 vildars 1
33524 vildaste 2
33525 vildmark 1
33526 vildmarken 2
33527 vildmarkens 1
33528 vilja 498
33529 viljan 22
33530 viljans 1
33531 viljekraft 1
33532 viljemässigt 1
33533 viljestark 1
33534 viljestarka 1
33535 vilka 267
33536 vilkas 10
33537 vilken 218
33538 vilket 608
33539 vill 1479
33540 village 1
33541 ville 81
33542 villervalla 1
33543 villig 8
33544 villiga 2
33545 villighet 2
33546 villigt 2
33547 villkor 85
33548 villkorande 1
33549 villkorar 1
33550 villkoren 30
33551 villkoret 1
33552 villkorliga 1
33553 villkorsuttryck 2
33554 villor 2
33555 villovägar 1
33556 villrådighet 1
33557 vilse 2
33558 vilsekommet 1
33559 vilseleda 2
33560 vilseledande 3
33561 vilseletts 1
33562 vilt 3
33563 vin 14
33564 vind 5
33565 vindar 2
33566 vinden 2
33567 vindfällen 1
33568 vindfällena 3
33569 vindlande 1
33570 vindruta 1
33571 vindskyffe 1
33572 vinet 3
33573 vingla 1
33574 vinkade 3
33575 vinkande 1
33576 vinkelräta 2
33577 vinklade 1
33578 vinklar 1
33579 vinkling 1
33580 vinna 11
33581 vinnande 1
33582 vinnare 1
33583 vinnarna 1
33584 vinnas 1
33585 vinner 4
33586 vinning 1
33587 vinodlingen 1
33588 vinproduktionen 1
33589 vinsektorn 1
33590 vinst 9
33591 vinsten 3
33592 vinster 17
33593 vinsterna 4
33594 vinstinriktade 2
33595 vinstintresse 2
33596 vinstintresset 2
33597 vinstjakt 1
33598 vinstmarginaler 1
33599 vinstsvag 1
33600 vinsttänkande 1
33601 vint 1
33602 vinter 1
33603 vintereftermiddag 1
33604 vintern 3
33605 vintertid 1
33606 vinthunds 1
33607 vinylfodral 1
33608 violer 1
33609 vippade 1
33610 vippen 1
33611 vira 1
33612 virka 1
33613 virkesförsäljning 1
33614 virkeslager 1
33615 virkeslagren 1
33616 virrigt 1
33617 virrvarr 1
33618 virtuellt 2
33619 virus 4
33620 virusbärare 1
33621 viruset 8
33622 virussjukdom 2
33623 virveln 2
33624 virvelvind 1
33625 virvlade 2
33626 virvlande 1
33627 vis 30
33628 visa 95
33629 visade 24
33630 visades 1
33631 visar 148
33632 visare 1
33633 visas 21
33634 visat 79
33635 visats 2
33636 visavi 2
33637 visdom 1
33638 vise 1
33639 visering 1
33640 viseringar 1
33641 viserings- 1
33642 vises 1
33643 viset 11
33644 vishet 1
33645 vishetens 1
33646 vision 17
33647 visionen 3
33648 visioner 9
33649 visiteras 1
33650 viskade 2
33651 viskades 1
33652 visningsformat 1
33653 vispgrädde 1
33654 viss 104
33655 vissa 378
33656 visselpipan 1
33657 visserligen 31
33658 visshet 3
33659 vissheten 1
33660 visslade 1
33661 visslande 1
33662 visst 32
33663 visste 45
33664 vistades 1
33665 vistas 4
33666 vistats 1
33667 vistelse 1
33668 vistelseort 1
33669 visualisera 1
33670 visuella 2
33671 visum 1
33672 vit 15
33673 vita 31
33674 vital 2
33675 vitala 3
33676 vitalisera 1
33677 vitaliseras 1
33678 vitalitet 1
33679 vitaliteten 1
33680 vitas 1
33681 vitaste 1
33682 vitblonda 1
33683 vitblänkande 1
33684 vitbok 34
33685 vitboken 44
33686 vitbokens 2
33687 vitbokssyndromet 1
33688 vitböcker 1
33689 vitböckerna 1
33690 vitglöd 1
33691 vitkalkade 1
33692 vitrinskåp 1
33693 vits 1
33694 vitt 11
33695 vittgående 1
33696 vittna 3
33697 vittnade 1
33698 vittnar 6
33699 vittnat 1
33700 vittne 3
33701 vittnen 1
33702 vittnesbördet 1
33703 vittnesförhör 1
33704 vittnet 1
33705 vittomfattande 4
33706 vittrande 1
33707 vittrar 1
33708 vitögat 1
33709 vivendi 2
33710 vokabulär 2
33711 volet 2
33712 voluntarism 2
33713 voluntaristiska 4
33714 volym 1
33715 volymen 2
33716 volymer 1
33717 von 23
33718 vore 82
33719 votering 1
33720 voteringssystemet 2
33721 votre 1
33722 votum 1
33723 vrak 6
33724 vrakdelarna 1
33725 vraket 3
33726 vrakets 1
33727 vrakgods 1
33728 vred 1
33729 vrede 3
33730 vreden 1
33731 vredgat 1
33732 vredgats 1
33733 vrida 3
33734 vrider 1
33735 vrist 1
33736 vräkte 1
33737 vräkts 2
33738 vrålade 2
33739 vrålande 1
33740 vulkanen 1
33741 vunnen 1
33742 vunnet 2
33743 vunnit 7
33744 vuxit 3
33745 vuxna 6
33746 vy 1
33747 vyer 5
33748 vykort 1
33749 vyn 2
33750 väcka 9
33751 väckarklocka 2
33752 väcker 11
33753 väcks 2
33754 väckt 4
33755 väckte 4
33756 väcktes 4
33757 väckts 2
33758 väder 2
33759 väderkvarnar 1
33760 väders 1
33761 väderstreck 2
33762 vädja 6
33763 vädjan 9
33764 vädjanden 4
33765 vädjar 12
33766 vädjat 1
33767 vädret 3
33768 väg 118
33769 väg- 1
33770 väga 7
33771 vägar 29
33772 vägarna 9
33773 vägas 2
33774 vägbyggnad 1
33775 vägde 1
33776 vägen 68
33777 väger 4
33778 vägg 4
33779 väggar 1
33780 väggarna 6
33781 väggen 7
33782 vägkontroller 4
33783 vägkontrollerna 1
33784 vägleda 1
33785 vägledande 8
33786 vägledning 2
33787 väglett 3
33788 vägmärken 1
33789 vägnar 42
33790 vägnät 1
33791 vägra 10
33792 vägrade 6
33793 vägran 11
33794 vägrar 13
33795 vägras 1
33796 vägrat 6
33797 vägröjare 1
33798 vägskäl 1
33799 vägskälet 1
33800 vägsträckan 1
33801 vägsäkerhetens 1
33802 vägtrafikanter 1
33803 vägtrafikants 1
33804 vägtrafiken 1
33805 vägtrafiksäkerheten 1
33806 vägtransporter 1
33807 väktare 6
33808 väl 177
33809 välbalanserad 2
33810 välbalanserade 2
33811 välbefinnande 2
33812 välbehövligt 1
33813 välbekant 2
33814 välbekanta 1
33815 välbeställda 1
33816 väldig 8
33817 väldiga 6
33818 väldigt 68
33819 välformade 1
33820 välformat 1
33821 välfunna 1
33822 välfärd 14
33823 välfärden 4
33824 välfärdsmässiga 1
33825 välfärdsmålen 1
33826 välfärdsnivån 1
33827 välfärdspolitiken 1
33828 välfärdssamhälle 1
33829 välfärdsskillnader 1
33830 välfärdsstaten 3
33831 välfärdsvinster 1
33832 välförvaltad 1
33833 välgrundad 2
33834 välgrundade 1
33835 välgång 1
33836 välgörande 3
33837 välinformerad 1
33838 välja 40
33839 väljarbastioner 1
33840 väljare 9
33841 väljarkåren 2
33842 väljarna 9
33843 väljarnas 2
33844 väljas 3
33845 väljer 21
33846 väljs 2
33847 välklingande 1
33848 välkommen 9
33849 välkommet 10
33850 välkomna 39
33851 välkomnade 2
33852 välkomnande 1
33853 välkomnar 87
33854 välkomnas 6
33855 välkomnat 1
33856 välkomnats 1
33857 välkomsthälsning 1
33858 välkvalificerade 1
33859 välkända 6
33860 välkänt 5
33861 vällde 1
33862 väller 1
33863 välmenande 1
33864 välment 1
33865 välmenta 2
33866 välmotiverad 1
33867 välmående 7
33868 välsignad 1
33869 välsignade 1
33870 välsignelse 1
33871 välsignelser 1
33872 välskött 1
33873 välstrukturerad 1
33874 välstånd 22
33875 välståndet 1
33876 välståndets 1
33877 välståndsnivå 1
33878 välståndsutvecklingen 1
33879 välta 1
33880 vältalig 1
33881 vältaligt 2
33882 vältra 1
33883 välutbildad 2
33884 välutbildade 1
33885 välutvecklad 1
33886 välutvecklade 1
33887 välvde 1
33888 vämjelse 1
33889 vän 23
33890 vända 23
33891 vändas 1
33892 vände 17
33893 vänder 16
33894 vändning 5
33895 vändningen 2
33896 vändpunkt 10
33897 vänja 1
33898 vänlig 4
33899 vänliga 3
33900 vänligen 4
33901 vänlighet 1
33902 vänligt 3
33903 vänner 26
33904 vännerna 1
33905 vänorter 1
33906 vänskap 5
33907 vänskapliga 1
33908 vänskapligt 1
33909 vänskapsband 1
33910 vänster 24
33911 vänsterbetänkande 1
33912 vänsterkritiker 1
33913 vänstern 16
33914 vänsterns 2
33915 vänsterregeringar 2
33916 vänsterregeringarna 1
33917 vänsterregeringens 1
33918 vänstra 3
33919 vänt 4
33920 vänta 43
33921 väntad 1
33922 väntade 18
33923 väntan 15
33924 väntar 47
33925 väntas 1
33926 väntat 11
33927 vänts 1
33928 väpnad 2
33929 väpnade 12
33930 värd 13
33931 värda 8
33932 värde 33
33933 värdedata 1
33934 värdefull 7
33935 värdefulla 10
33936 värdefullt 5
33937 värdegemenskap 5
33938 värdegrund 1
33939 värdelös 2
33940 värdelösa 2
33941 värdemässigt 1
33942 värden 41
33943 värdena 8
33944 värdenamn 2
33945 värdepapper 6
33946 värdepappersfonder 1
33947 värdepappersfondernas 1
33948 värdepappersmarknaden 1
33949 värdepappersområdet 2
33950 värdera 2
33951 värderade 7
33952 värderar 2
33953 värderas 5
33954 värdering 3
33955 värderingar 36
33956 värderingarna 4
33957 värderingarnas 1
33958 värdestegring 1
33959 värdesystem 1
33960 värdesätta 1
33961 värdesätter 1
33962 värdet 14
33963 värdeökningen 1
33964 värdig 3
33965 värdighet 14
33966 värdigheten 2
33967 värdigt 4
33968 värdinna 1
33969 värdinnorna 1
33970 värdlandet 1
33971 värdmedlemsstatens 1
33972 värja 1
33973 värjer 1
33974 värkande 1
33975 värkar 1
33976 värld 30
33977 världar 3
33978 världen 160
33979 världens 39
33980 världsbefolkningen 1
33981 världsbild 1
33982 världsdel 6
33983 världsdelar 2
33984 världsdelen 3
33985 världsekonomin 7
33986 världsfinansens 1
33987 världsfrågorna 1
33988 världsfrånvända 1
33989 världshandel 2
33990 världshandeln 3
33991 världshandelsförhandlingar 1
33992 världskonferens 2
33993 världskrig 1
33994 världskriget 5
33995 världskrigets 3
33996 världsledande 1
33997 världsliga 1
33998 världsmakts 1
33999 världsmarknaden 4
34000 världsmarknaderna 1
34001 världsmedborgare 1
34002 världsmodell 1
34003 världsnivå 1
34004 världsomspännande 7
34005 världsordning 3
34006 världsordningen 2
34007 världsregering 1
34008 världsriken 1
34009 världssamfundet 7
34010 världssamfundets 1
34011 världsstandard 1
34012 världsstyre 1
34013 världsuppfattning 1
34014 världsvana 1
34015 världsvattenforum 1
34016 världsövergripande 1
34017 värmas 1
34018 värmde 3
34019 värme 3
34020 värmen 2
34021 värmepannan 1
34022 värmt 1
34023 värna 9
34024 värnar 6
34025 värre 15
34026 värst 3
34027 värsta 23
34028 värt 14
34029 värv 2
34030 värvas 1
34031 väsande 1
34032 väsen 3
34033 väsendet 1
34034 väsentlig 17
34035 väsentliga 19
34036 väsentligen 2
34037 väsentligheterna 1
34038 väsentligt 23
34039 väska 3
34040 väskan 2
34041 väskorna 1
34042 väst 3
34043 västafrikanska 1
34044 väster 2
34045 västerländsk 1
34046 västerländska 1
34047 västern 1
34048 västerut 1
34049 västeuropeiska 1
34050 västkusten 1
34051 västliga 1
34052 västländerna 3
34053 västländernas 1
34054 västra 7
34055 västvärlden 2
34056 väv 1
34057 vävnad 3
34058 vävnaden 1
34059 vävnader 1
34060 vävt 1
34061 växa 11
34062 växande 15
34063 växandets 1
34064 växelkontor 1
34065 växelkursen 1
34066 växelkurser 1
34067 växelkurserna 1
34068 växelkurspolitiken 1
34069 växelkursutvecklingen 1
34070 växelspel 1
34071 växelverkan 2
34072 växer 17
34073 växla 2
34074 växlande 1
34075 växlar 2
34076 växlas 1
34077 växlat 2
34078 växling 1
34079 växlingarna 2
34080 växtarter 1
34081 växte 6
34082 växter 3
34083 växtfrämjande 1
34084 växthuseffekt 1
34085 växthuseffekten 5
34086 växthusgaser 4
34087 växthusgaserna 2
34088 växtliv 2
34089 växtskydd 2
34090 växtskyddsproblem 1
34091 våg 2
34092 våga 3
34093 vågade 4
34094 vågar 13
34095 vågat 3
34096 vågen 1
34097 vågiga 1
34098 våglängd 1
34099 vågor 1
34100 vågorna 1
34101 vågrät 2
34102 vågskålen 1
34103 våld 12
34104 våldet 13
34105 våldets 2
34106 våldsam 4
34107 våldsamhet 1
34108 våldsamma 6
34109 våldsamt 3
34110 våldsbenägen 1
34111 våldsdemonstrationer 1
34112 våldsdåd 1
34113 våldsdåden 1
34114 våldshandlingar 2
34115 våldskultur 1
34116 våldsuttryck 1
34117 våldta 1
34118 våldtagen 1
34119 våldtagits 1
34120 våldtas 2
34121 våldtogs 1
34122 våldtäkt 2
34123 våldtäkter 1
34124 våldtäkterna 1
34125 vållade 1
34126 vållar 3
34127 våning 2
34128 våningar 1
34129 våningen 3
34130 vår 520
34131 våra 483
34132 vård 3
34133 vårda 1
34134 vårdad 1
34135 vårdade 1
34136 vårdar 3
34137 vårdcentraler 1
34138 vården 1
34139 vårdslös 1
34140 vårdslöshet 2
34141 våren 3
34142 vårens 1
34143 vårt 308
34144 våta 1
34145 våtare 1
34146 våtmarksområden 1
34147 våtområden 1
34148 vått 1
34149 vördnad 3
34150 vördnadsvärda 1
34151 walesare 1
34152 walesiska 1
34153 wallonska 1
34154 webben 1
34155 webbläsare 1
34156 webbläsaren 2
34157 webbplats 2
34158 webbsida 4
34159 webbsidan 1
34160 webbsidans 1
34161 webbsidor 1
34162 webbsidorna 1
34163 weitergeführt 1
34164 welfare 1
34165 werden 1
34166 whisky 6
34167 with 3
34168 within 1
34169 worst 1
34170 yawlen 1
34171 yen 1
34172 ylle 1
34173 yllesjalar 1
34174 yngelperioder 1
34175 yngre 3
34176 yngsta 1
34177 ynkliga 1
34178 ynkligt 1
34179 yppas 1
34180 ypperligt 2
34181 yppig 1
34182 yrka 7
34183 yrkande 6
34184 yrkanden 2
34185 yrkandet 2
34186 yrkar 8
34187 yrkat 1
34188 yrken 4
34189 yrkes- 1
34190 yrkesaktivas 1
34191 yrkesarbetande 2
34192 yrkesetik 1
34193 yrkesfiskarna 3
34194 yrkesfiskarnas 2
34195 yrkesgrupper 3
34196 yrkesjurister 1
34197 yrkeskarriärer 1
34198 yrkeskunnande 1
34199 yrkeskvalifikationer 2
34200 yrkeslivet 4
34201 yrkeslivets 1
34202 yrkesman 1
34203 yrkesmässig 1
34204 yrkesmässiga 2
34205 yrkesmässigt 1
34206 yrkesområdet 1
34207 yrkesprofil 1
34208 yrkestrafik 1
34209 yrkesutbildning 10
34210 yrkesutbildningen 2
34211 yrkesutbildningsåtgärder 1
34212 yrkesval 1
34213 yrkesverksamheter 1
34214 yrkesverksamma 7
34215 yrsel 1
34216 yt- 2
34217 yta 6
34218 ytan 4
34219 ytlig 1
34220 ytliga 1
34221 ytlighet 1
34222 ytligt 1
34223 ytorna 1
34224 ytskeendet 1
34225 ytterdörren 3
34226 ytterkläder 1
34227 ytterligare 182
34228 ytterligheten 3
34229 ytterligheter 1
34230 ytterlighetsåtgärder 1
34231 ytterligt 3
34232 ytterområde 1
34233 ytterområden 2
34234 ytterskrovet 1
34235 ytterst 61
34236 yttersta 34
34237 yttertrappan 1
34238 yttervärlden 2
34239 yttra 11
34240 yttrande 41
34241 yttrandefrihet 3
34242 yttranden 5
34243 yttrandet 13
34244 yttrar 2
34245 yttrat 1
34246 yttrats 3
34247 yttre 26
34248 ytvatten 9
34249 ytvattenstatus 2
34250 ytvattnen 1
34251 ytvattnens 1
34252 ytvattnet 8
34253 yviga 1
34254 yxa 1
34255 zero 1
34256 zigenare 3
34257 zigenarflyktingar 1
34258 zigenarna 1
34259 zigenska 1
34260 zon 2
34261 zoner 1
34262 zoners 1
34263 zonindelningen 1
34264 zu 9
34265 § 1
34266 ­ 1
34267 ­företräds 1
34268 ­inom 1
34269 º 1
34270 ¿ 1
34271 Álvaro 2
34272 Äldre 1
34273 Ämnar 1
34274 Ämnet 1
34275 Än 10
34276 Ända 6
34277 Ändra 4
34278 Ändras 1
34279 Ändringar 1
34280 Ändringsförslag 35
34281 Ändringsförslagen 11
34282 Ändå 24
34283 Ännu 11
34284 Äntligen 4
34285 Är 71
34286 Ärade 33
34287 Ärendet 1
34288 Ärkebiskopen 1
34289 Ärret 2
34290 Ät 1
34291 Även 122
34292 Å 65
34293 Åhå 1
34294 Åklagaren 1
34295 Ånyo 1
34296 År 12
34297 Året 1
34298 Årligen 1
34299 Årligt 1
34300 Åsikt 2
34301 Åt 1
34302 Åtagandet 1
34303 Åtal 1
34304 Återetableringslagen 1
34305 Återigen 2
34306 Återinrättandet 1
34307 Återspeglas 1
34308 Återstående 1
34309 Återstår 2
34310 Återupptagande 6
34311 Återvinningskraven 1
34312 Åtgärd 1
34313 Åtgärder 10
34314 Åtgärderna 2
34315 Åtgärdernas 1
34316 Åtminstone 2
34317 Åtta 1
34318 Émilie 1
34319 Ésclope 1
34320 Île-de-France 1
34321 ÖVP 9
34322 Ödet 1
34323 Ögonblicket 3
34324 Ögonen 1
34325 Öh 1
34326 Ökad 1
34327 Ön 1
34328 Önskar 1
34329 Önskemålet 1
34330 Öppenhet 2
34331 Öppna 1
34332 Öppnande 1
34333 Öst- 1
34334 Österrike 99
34335 Österrikes 14
34336 Österrikiska 11
34337 Östersjöländerna 1
34338 Östersjön 5
34339 Östersjöområdet 1
34340 Östersjöregionens 1
34341 Östeuropa 18
34342 Östeuropas 1
34343 Östtimor 8
34344 Östturkestan 1
34345 Östtyskland 4
34346 Över 6
34347 Överallt 1
34348 Överfisket 1
34349 Övergrepp 1
34350 Övergreppen 1
34351 Överproduktionen 1
34352 Överst 1
34353 Överste 2
34354 Översvämningar 1
34355 Översvämningarna 1
34356 Överväger 1
34357 Övriga 2
34358 à 1
34359 äcklar 1
34360 ädelstenar 2
34361 ädelt 2
34362 ädla 1
34363 äga 71
34364 ägandeform 1
34365 ägandeförhållanden 2
34366 äganderätten 1
34367 ägandet 1
34368 ägaransvaret 1
34369 ägare 10
34370 ägaren 8
34371 ägares 1
34372 ägarna 2
34373 ägarnas 1
34374 ägas 1
34375 ägde 13
34376 äger 33
34377 ägg 2
34378 ägna 23
34379 ägnad 1
34380 ägnade 7
34381 ägnar 29
34382 ägnas 4
34383 ägnat 9
34384 ägnats 1
34385 ägodelar 3
34386 ägt 15
34387 äkta 9
34388 äktenskap 2
34389 äktenskapsmål 1
34390 äldre 43
34391 äldreomsorg 1
34392 äldreomsorgen 1
34393 äldres 4
34394 äldsta 4
34395 älska 5
34396 älskade 8
34397 älskar 6
34398 älskare 1
34399 älskvärd 1
34400 älskvärda 2
34401 älskvärdhet 1
34402 älvar 1
34403 ämbete 6
34404 ämbetsmannalagen 1
34405 ämbetsmännen 1
34406 ämbetsrum 1
34407 ämna 1
34408 ämnade 3
34409 ämnar 9
34410 ämne 42
34411 ämnen 62
34412 ämnena 9
34413 ämnesområde 2
34414 ämnesområdena 1
34415 ämnesprioriteringarna 1
34416 ämnet 15
34417 ämnets 1
34418 än 606
34419 ända 25
34420 ändamål 12
34421 ändamålen 1
34422 ändamålet 12
34423 ändamålsenlig 5
34424 ändamålsenliga 5
34425 ändamålsenligheten 2
34426 ändamålsenligt 4
34427 ändarna 1
34428 ände 5
34429 änden 2
34430 ändlös 2
34431 ändlösa 5
34432 ändock 1
34433 ändpunkter 1
34434 ändra 76
34435 ändrad 3
34436 ändrade 6
34437 ändrades 1
34438 ändrar 11
34439 ändras 26
34440 ändrat 9
34441 ändrats 9
34442 ändring 61
34443 ändringar 69
34444 ändringarna 13
34445 ändringen 11
34446 ändringsakter 1
34447 ändringsdirektiv 1
34448 ändringsförlag 1
34449 ändringsförslag 431
34450 ändringsförslagen 81
34451 ändringsförslaget 21
34452 ändringsförslagets 1
34453 ändå 161
34454 ängarna 2
34455 ängel 1
34456 ängels 1
34457 ängen 1
34458 ängslan 2
34459 ängsliga 2
34460 ängsligt 3
34461 änka 1
34462 ännu 241
34463 äntligen 67
34464 äntrade 1
34465 är 8224
34466 ära 1
34467 ärade 116
34468 äran 10
34469 ärende 36
34470 ärenden 8
34471 ärendena 6
34472 ärendet 20
34473 ärendets 1
34474 ärkefiende 1
34475 ärlig 4
34476 ärliga 6
34477 ärlighet 1
34478 ärligt 11
34479 ärmarna 1
34480 ärmen 1
34481 äro 1
34482 ärofylld 1
34483 ärr 2
34484 ärrbildning 1
34485 ärret 1
34486 ärvt 1
34487 ät 1
34488 äta 18
34489 ätas 1
34490 äter 7
34491 ätit 2
34492 ättning 1
34493 även 811
34494 äventyr 2
34495 äventyra 11
34496 äventyrades 1
34497 äventyrar 14
34498 äventyrare 1
34499 äventyras 4
34500 å 92
34501 åberopa 4
34502 åberopar 1
34503 åberopas 1
34504 ådra 1
34505 ådrog 1
34506 ådror 2
34507 ådrorna 1
34508 åh 1
34509 åhörare 1
34510 åhörarläktaren 3
34511 åhörarläktarna 1
34512 åhört 1
34513 åka 8
34514 åker 2
34515 åkerier 1
34516 åkern 1
34517 åklagare 20
34518 åklagaren 8
34519 åklagares 1
34520 åklagarmyndighet 9
34521 åklagarmyndigheten 4
34522 åklagarmyndigheter 1
34523 åklagarna 1
34524 åklagarämbete 1
34525 åkommor 1
34526 åkte 2
34527 ål 2
34528 ålagd 2
34529 ålagda 2
34530 ålagts 2
34531 ålder 16
34532 ålderdomen 1
34533 ålderdomlig 1
34534 ålderdomshem 2
34535 åldern 2
34536 ålders 1
34537 ålderspensionen 1
34538 ålderstigen 1
34539 ålderstigna 1
34540 åldersökning 1
34541 åldrade 1
34542 åldrande 5
34543 åldrandet 1
34544 åldras 1
34545 åldrats 1
34546 åldringar 1
34547 åligga 3
34548 åligger 7
34549 ålägga 5
34550 ålägganden 1
34551 åläggandet 1
34552 åläggas 1
34553 ålägger 6
34554 åläggs 1
34555 ån 1
34556 ångare 2
34557 ångat 1
34558 ångbåtar 1
34559 ånger 1
34560 ångestfyllda 1
34561 ångestfyllt 1
34562 ånglok 1
34563 ångorna 1
34564 ångpanna 1
34565 ångrade 1
34566 ångvälten 1
34567 ånyo 3
34568 år 580
34569 år- 1
34570 åra 1
34571 åratal 9
34572 åren 126
34573 årens 13
34574 året 88
34575 årets 7
34576 århundrade 7
34577 århundraden 4
34578 århundradet 13
34579 århundradets 1
34580 årlig 6
34581 årliga 35
34582 årligen 14
34583 årligt 2
34584 års 42
34585 årsbeloppet 1
34586 årsberättelser 1
34587 årsrapport 3
34588 årsrapporten 2
34589 årsrapporter 1
34590 årstiden 1
34591 årsungar 2
34592 årsvis 1
34593 årtal 1
34594 årtionde 1
34595 årtionden 4
34596 årtiondena 1
34597 årtiondet 1
34598 årtusende 2
34599 årtusendena 1
34600 årtusendeskiftet 1
34601 årtusendet 1
34602 årtusendets 1
34603 åsamkar 1
34604 åsamkas 1
34605 åsamkat 4
34606 åsatt 1
34607 åsidosatte 1
34608 åsidosattes 2
34609 åsidosätta 3
34610 åsidosättande 2
34611 åsidosätter 3
34612 åsikt 74
34613 åsikten 8
34614 åsikter 37
34615 åsikterna 9
34616 åsiktsförbrytelser 1
34617 åsiktsförklaring 1
34618 åsiktsskillnad 1
34619 åsiktsskillnader 2
34620 åsiktsutbyten 1
34621 åskådarbalkongen 1
34622 åskådare 3
34623 åskådaren 1
34624 åskådliggjordes 1
34625 åskådning 1
34626 åsna 1
34627 åsnorna 1
34628 åstad 1
34629 åstadkom 2
34630 åstadkomma 39
34631 åstadkommas 3
34632 åstadkommer 7
34633 åstadkommit 6
34634 åstadkommits 3
34635 åstadkoms 1
34636 åsyftade 5
34637 åsyftar 5
34638 åsyftas 4
34639 åsynen 1
34640 åt 289
34641 åta 6
34642 åtagande 28
34643 åtagande- 1
34644 åtaganden 40
34645 åtagandena 4
34646 åtagandet 6
34647 åtagandetakt 1
34648 åtagit 10
34649 åtal 8
34650 åtala 3
34651 åtalade 2
34652 åtalas 4
34653 åtalsfasen 1
34654 åtalspunkter 3
34655 åtalspunkterna 3
34656 åtanke 8
34657 åtar 5
34658 åter 64
34659 återanpassa 1
34660 återanpassning 2
34661 återanställningsprocesserna 1
34662 återanvända 2
34663 återanvändas 1
34664 återanvändbara 1
34665 återanvändning 9
34666 återanvändningen 1
34667 återanvändnings- 1
34668 återanvändningsbart 1
34669 återanvändningsnivåer 1
34670 återanvänt 1
34671 återbetala 2
34672 återbetalats 1
34673 återbetalning 2
34674 återerövra 1
34675 återerövrande 1
34676 återerövring 1
34677 återetableringslag 1
34678 återfaller 1
34679 återfick 1
34680 återfinnas 2
34681 återfinner 2
34682 återfinns 6
34683 återfunna 1
34684 återfunnen 1
34685 återfå 1
34686 återfår 1
34687 återföras 2
34688 återfördela 1
34689 återfördes 1
34690 återförena 2
34691 återförenat 1
34692 återförening 1
34693 återföringen 1
34694 återförs 1
34695 återförts 1
34696 återförvisa 1
34697 återförvisas 3
34698 återförvisning 1
34699 återförvisningen 1
34700 återförvärva 1
34701 återgav 2
34702 återgavs 2
34703 återge 8
34704 återger 2
34705 återges 2
34706 återgett 1
34707 återgick 1
34708 återgivande 1
34709 återgivning 1
34710 återgå 2
34711 återgång 1
34712 återgår 1
34713 återgått 1
34714 återhämta 2
34715 återhämtning 9
34716 återhämtningen 4
34717 återhämtningsnivåer 1
34718 återhämtningsprogram 1
34719 återhållen 1
34720 återhållsam 1
34721 återhållsamhet 1
34722 återhållsamma 4
34723 återigen 50
34724 återinför 2
34725 återinföra 2
34726 återinförande 1
34727 återinförs 1
34728 återinresa 1
34729 återintagande 1
34730 återintegrering 1
34731 återintegreringsprogram 1
34732 återkalla 2
34733 återkallad 1
34734 återknyta 2
34735 återkom 1
34736 återkomma 6
34737 återkommande 5
34738 återkommer 6
34739 återkommit 1
34740 återkomst 1
34741 återkomsten 1
34742 återkräva 2
34743 återkrävas 1
34744 återlämna 3
34745 åternationalisera 3
34746 åternationaliseras 1
34747 åternationalisering 7
34748 åternationaliseringen 1
34749 återsamla 1
34750 återskapa 7
34751 återspegla 3
34752 återspeglar 6
34753 återspeglas 4
34754 återspegling 1
34755 återstod 1
34756 återställa 25
34757 återställande 4
34758 återställandet 2
34759 återställas 1
34760 återställer 1
34761 återställs 1
34762 återstående 3
34763 återstår 27
34764 återsända 1
34765 återsänds 1
34766 återta 2
34767 återtagande 4
34768 återtagandet 3
34769 återtar 1
34770 återtas 1
34771 återtog 1
34772 återuppbygga 2
34773 återuppbyggandet 5
34774 återuppbyggnad 8
34775 återuppbyggnaden 12
34776 återuppbyggnader 1
34777 återuppbyggnadsarbete 1
34778 återuppbyggnadsarbetena 1
34779 återuppbyggnadsfas 1
34780 återuppbyggnadsorgan 1
34781 återuppbyggnadsprogram 2
34782 återuppbyggnadsprogrammet 1
34783 återuppbyggt 1
34784 återuppfinna 1
34785 återuppliva 1
34786 återupplivande 1
34787 återupplivandet 1
34788 återupprepa 1
34789 återupprepas 3
34790 återupprätta 13
34791 återupprättandet 1
34792 återupprättar 2
34793 återupprättas 2
34794 återuppstå 1
34795 återuppståndelse 1
34796 återuppstår 1
34797 återuppstått 1
34798 återuppta 3
34799 återupptagande 1
34800 återupptagandet 2
34801 återupptagen 5
34802 återupptagits 1
34803 återupptagna 2
34804 återupptar 3
34805 återupptas 3
34806 återupptogs 13
34807 återupptäcka 1
34808 återuppvaknandet 1
34809 återverkan 1
34810 återverkningar 1
34811 återvinna 16
34812 återvinnande 2
34813 återvinnas 7
34814 återvinner 3
34815 återvinning 22
34816 återvinningen 6
34817 återvinningsbart 1
34818 återvinningsföretag 1
34819 återvinningsgrad 1
34820 återvinningsindustrin 1
34821 återvinningskostnaderna 2
34822 återvinningskravet 1
34823 återvinningsmodell 1
34824 återvinningsmonopol 1
34825 återvinningsmål 2
34826 återvinningsmålet 1
34827 återvinningsprocessen 1
34828 återvinningssektor 1
34829 återvinningssektorn 1
34830 återvinningssystem 1
34831 återvinningsverksamheten 1
34832 återvinningsvänliga 1
34833 återvinns 2
34834 återvunna 1
34835 återvunnet 1
34836 återvända 7
34837 återvände 2
34838 återvänder 4
34839 återvändsgränd 2
34840 återvänt 2
34841 åtfölja 5
34842 åtföljande 4
34843 åtföljas 8
34844 åtföljde 1
34845 åtföljdes 1
34846 åtföljer 1
34847 åtföljs 6
34848 åtföljt 1
34849 åtföljts 1
34850 åtgärd 47
34851 åtgärda 2
34852 åtgärdar 2
34853 åtgärdas 5
34854 åtgärden 8
34855 åtgärdens 1
34856 åtgärder 446
34857 åtgärderna 37
34858 åtgärds 1
34859 åtgärdsgrupper 1
34860 åtgärdsgrupperna 1
34861 åtgärdslista 2
34862 åtgärdsområden 1
34863 åtgärdspaket 7
34864 åtgärdspaketet 1
34865 åtgärdsplan 4
34866 åtgärdsplanen 1
34867 åtgärdsplanerna 1
34868 åtgärdsprogram 9
34869 åtgärdsprogrammen 2
34870 åtgärdsprogrammet 1
34871 åtgärdspunkter 1
34872 åtgärdsrelaterade 1
34873 åthävor 1
34874 åtkomlig 1
34875 åtlydd 1
34876 åtminstone 94
34877 åtnjuta 6
34878 åtnjutande 1
34879 åtnjuter 3
34880 åtnjöt 1
34881 åtog 3
34882 åtrådd 1
34883 åtrådde 2
34884 åtrår 1
34885 åtråvärdhet 1
34886 åtskilda 1
34887 åtskilja 1
34888 åtskillig 1
34889 åtskilliga 3
34890 åtskilligt 1
34891 åtskillnad 5
34892 åtstramning 4
34893 åtstramningar 2
34894 åtta 14
34895 åttasidiga 1
34896 åttatiden 1
34897 åttonde 2
34898 åvilar 3
34899 ö 6
34900 öar 2
34901 öarna 12
34902 öarnas 1
34903 öbo 1
34904 öbor 1
34905 öde 31
34906 ödelade 2
34907 ödelagd 1
34908 ödelagda 2
34909 ödelägga 1
34910 ödeläggande 1
34911 ödeläggelse 2
34912 ödeläggelsen 1
34913 ödeläggs 1
34914 ödemark 2
34915 ödemarken 1
34916 öden 1
34917 ödesbestämda 1
34918 ödesbestämt 1
34919 ödesdiger 1
34920 ödesdigert 2
34921 ödesdigra 4
34922 ödesgemenskap 3
34923 ödesmättade 1
34924 ödet 1
34925 ödslig 1
34926 öga 8
34927 ögat 4
34928 ögla 1
34929 ögon 46
34930 ögonblick 55
34931 ögonblicken 2
34932 ögonblicket 22
34933 ögonblickligen 1
34934 ögonen 14
34935 ögonfärg 1
34936 ögontjänarna 1
34937 ögonvitor 1
34938 öka 98
34939 ökad 68
34940 ökade 27
34941 ökades 1
34942 ökande 14
34943 ökar 50
34944 ökas 7
34945 ökat 39
34946 öken 1
34947 ökenområden 1
34948 ökenområdet 1
34949 ökenspridningen 1
34950 ökenutbredning 2
34951 ökenutbredningen 1
34952 öknar 1
34953 öknen 1
34954 ökning 32
34955 ökningen 8
34956 ökningseffekt 1
34957 ökningsprincipen 1
34958 öl 5
34959 ölflaskorna 1
34960 ölkrus 1
34961 ölsort 1
34962 öm 1
34963 ömma 1
34964 ömmande 1
34965 ömsesidig 10
34966 ömsesidiga 5
34967 ömsesidighet 1
34968 ömsesidigt 9
34969 ömtåliga 3
34970 ömtålighet 1
34971 ömänniskor 1
34972 ön 21
34973 öns 6
34974 önska 21
34975 önskad 3
34976 önskade 8
34977 önskan 35
34978 önskar 56
34979 önskas 1
34980 önskat 5
34981 önskelista 1
34982 önskelistan 1
34983 önskelistor 1
34984 önskemål 16
34985 önskemålen 2
34986 önsketänkandet 1
34987 önskning 1
34988 önskningar 6
34989 önskvärd 6
34990 önskvärda 3
34991 önskvärt 18
34992 öområden 2
34993 öområdena 1
34994 öppen 35
34995 öppenhet 89
34996 öppenheten 17
34997 öppenhetens 1
34998 öppenhets- 1
34999 öppenhetslag 1
35000 öppenhetslagstiftning 1
35001 öppet 36
35002 öppettider 1
35003 öppna 45
35004 öppnad 1
35005 öppnade 11
35006 öppnades 3
35007 öppnandet 1
35008 öppnar 20
35009 öppnare 3
35010 öppnas 7
35011 öppnat 2
35012 öppnats 2
35013 öppning 4
35014 öppningar 3
35015 öppningsanförande 1
35016 öppningsanförandet 1
35017 öppningserbjudande 1
35018 öppningshögtid 1
35019 öra 5
35020 öre 2
35021 öregion 1
35022 öregioner 5
35023 öregionerna 9
35024 örlogsmannen 1
35025 örngott 1
35026 örnnäsa 1
35027 öron 6
35028 öronbedövande 2
35029 öronen 3
35030 öronmärka 1
35031 öronmärkta 1
35032 ösa 1
35033 ösamhällen 1
35034 öst 4
35035 öst- 2
35036 östaterna 2
35037 östblocket 1
35038 öste 2
35039 öster 4
35040 österländska 1
35041 östern 2
35042 österrikare 3
35043 österrikarens 1
35044 österrikares 1
35045 österrikarna 5
35046 österrikisk 5
35047 österrikiska 56
35048 österrikiske 2
35049 österrikiskt 1
35050 österut 2
35051 östeuropeiska 5
35052 östländerna 2
35053 östländernas 1
35054 östra 9
35055 östrepublikerna 1
35056 östutvidgningen 2
35057 öva 1
35058 övat 1
35059 över 675
35060 överallt 23
35061 överarmen 1
35062 överbefolkade 1
35063 överbefälhavare 1
35064 överbelasta 1
35065 överbelastad 3
35066 överbemanning 1
35067 överblick 1
35068 överblicka 1
35069 överblivna 1
35070 överbord 2
35071 överbringa 1
35072 överbrygga 4
35073 överbryggas 1
35074 överbud 4
35075 övercentralisering 1
35076 överdimensionerad 1
35077 överdrift 2
35078 överdrifter 1
35079 överdriva 1
35080 överdrivas 1
35081 överdriven 12
35082 överdriver 3
35083 överdrivet 8
35084 överdrivna 5
35085 överdåd 1
35086 överdådiga 1
35087 överens 107
35088 överenskommelse 38
35089 överenskommelsen 6
35090 överenskommelser 5
35091 överenskommelserna 1
35092 överenskommen 1
35093 överenskommet 1
35094 överenskommits 2
35095 överenskomna 5
35096 överensstämde 1
35097 överensstämma 6
35098 överensstämmande 3
35099 överensstämmelse 19
35100 överensstämmer 21
35101 överexploatering 1
35102 överfall 3
35103 överfiske 2
35104 överfiskning 1
35105 överflyttas 1
35106 överflyttning 2
35107 överflödig 2
35108 överflödigt 3
35109 överfulla 1
35110 överföll 3
35111 överför 5
35112 överföra 9
35113 överförande 1
35114 överföras 6
35115 överförda 1
35116 överföring 20
35117 överföringar 2
35118 överföringarna 1
35119 överföringen 5
35120 överförs 6
35121 överförts 1
35122 övergav 1
35123 överge 4
35124 överger 6
35125 överges 5
35126 övergick 1
35127 övergiven 1
35128 övergivenhet 1
35129 övergivit 1
35130 övergivits 3
35131 övergivna 5
35132 övergrepp 2
35133 övergripande 32
35134 övergå 3
35135 övergång 6
35136 övergången 8
35137 övergångs- 1
35138 övergångsbestämmelser 3
35139 övergångsbestämmelserna 1
35140 övergångsfas 1
35141 övergångsperiod 6
35142 övergångsperioden 5
35143 övergångsperiodens 1
35144 övergångsperioder 1
35145 övergångssystemet 2
35146 övergångsår 1
35147 övergår 6
35148 övergått 1
35149 övergödd 1
35150 överhanden 1
35151 överhuvud 2
35152 överhuvudtaget 8
35153 överhängande 2
35154 överhöghet 3
35155 överilat 2
35156 överinseende 2
35157 överkastet 1
35158 överklaga 2
35159 överklagande 2
35160 överklagandeförfarande 1
35161 överklaganden 2
35162 överklagar 1
35163 överklagat 1
35164 överkomliga 3
35165 överkomligt 1
35166 överkomma 1
35167 överkommit 1
35168 överkommits 1
35169 överkörd 1
35170 överlade 2
35171 överlagda 1
35172 överlagt 1
35173 överlappar 3
35174 överlappning 2
35175 överlappningar 1
35176 överledas 1
35177 överledning 1
35178 överledningar 1
35179 överledningarna 1
35180 överledningen 4
35181 överleva 11
35182 överlevandet 1
35183 överlevde 3
35184 överlever 3
35185 överlevnad 3
35186 överlevt 2
35187 överläggningar 7
35188 överläggningarna 2
35189 överlägsen 1
35190 överlägsenhet 2
35191 överlägsenheten 1
35192 överlämna 8
35193 överlämnad 1
35194 överlämnade 3
35195 överlämnades 3
35196 överlämnande 1
35197 överlämnandet 2
35198 överlämnar 15
35199 överlämnas 5
35200 överlämnat 4
35201 överlämnats 6
35202 överlåta 9
35203 överlåtandet 1
35204 överlåtas 1
35205 överlåtbara 4
35206 överlåtelse 1
35207 överlåtelser 1
35208 överlåter 1
35209 överlåtit 1
35210 överlåtits 1
35211 överlåts 2
35212 övermaskinist 1
35213 övermekaniserade 1
35214 övermodigt 1
35215 övermorgon 5
35216 övermänsklig 1
35217 övernationell 4
35218 övernationella 2
35219 övernitiska 1
35220 övernog 1
35221 överordnad 1
35222 överordnade 1
35223 överpriser 1
35224 överraskad 2
35225 överraskade 1
35226 överraskande 5
35227 överraskning 6
35228 överregionala 1
35229 överreglerande 1
35230 överreglerat 1
35231 överreglering 1
35232 överrock 2
35233 överrocken 2
35234 överrumplad 1
35235 överrumplat 1
35236 överräckande 1
35237 överrätten 1
35238 överrösta 1
35239 översatta 1
35240 översatte 1
35241 översattes 2
35242 översatts 1
35243 överseende 1
35244 översida 1
35245 översikt 6
35246 översikten 8
35247 översikter 1
35248 översiktsplan 1
35249 överskott 6
35250 överskottet 2
35251 överskottskapacitet 1
35252 överskridas 1
35253 överskrider 4
35254 överskridit 1
35255 överskridits 1
35256 överskrids 3
35257 överskriften 3
35258 överskugga 2
35259 överskuggar 1
35260 överskådlig 5
35261 överspänd 2
35262 överst 2
35263 överstat 1
35264 överstaten 1
35265 överstatliga 1
35266 överstatlighet 4
35267 överstatligt 1
35268 överste 1
35269 översteg 1
35270 överstiga 1
35271 överstiger 5
35272 överstigit 1
35273 överståndet 1
35274 överståndna 1
35275 översvämmade 2
35276 översvämmades 1
35277 översvämmas 1
35278 översvämning 2
35279 översvämningar 11
35280 översvämningarna 9
35281 översvämningsbistånd 1
35282 översvämningsproblem 1
35283 översyn 8
35284 översynen 2
35285 översänd 1
35286 översända 1
35287 översändes 1
35288 översänds 1
35289 översätta 2
35290 översättarhus 1
35291 översättas 1
35292 översättning 1
35293 översättningar 4
35294 översättningarna 3
35295 översättningen 5
35296 översättningsarbeten 1
35297 översättningsfelen 1
35298 översättningsmisstag 1
35299 översättningsproblem 2
35300 översättningsproblemet 1
35301 översättningstjänst 1
35302 översättningstjänsten 2
35303 översållad 1
35304 överta 8
35305 övertag 2
35306 övertagande 1
35307 övertaganden 1
35308 övertagits 1
35309 övertala 1
35310 övertalade 1
35311 övertar 1
35312 övertid 1
35313 övertog 2
35314 övertoner 1
35315 övertramp 2
35316 överträdde 1
35317 överträdelse 3
35318 överträdelser 15
35319 överträdelserna 1
35320 överträds 2
35321 överträffa 1
35322 överträffar 1
35323 övertyga 17
35324 övertygad 50
35325 övertygade 18
35326 övertygande 15
35327 övertygar 1
35328 övertygat 4
35329 övertygelse 16
35330 övertygelsen 3
35331 övertygelsers 1
35332 övertänkta 1
35333 övervaka 18
35334 övervakade 1
35335 övervakar 2
35336 övervakas 7
35337 övervakat 1
35338 övervakning 19
35339 övervakningen 6
35340 övervakningscentra 2
35341 övervakningscentrer 1
35342 övervakningscentrum 4
35343 övervakningsformer 1
35344 övervakningsinstans 1
35345 övervakningssystem 1
35346 överviktig 1
35347 övervinna 10
35348 övervinnas 1
35349 övervinner 1
35350 övervinns 1
35351 övervunnits 1
35352 överväga 36
35353 övervägande 7
35354 överväganden 10
35355 övervägas 2
35356 övervägd 1
35357 övervägda 1
35358 övervägde 1
35359 överväger 12
35360 övervägs 1
35361 övervägt 2
35362 överväldigande 9
35363 övervältra 1
35364 övervåningen 1
35365 överösa 1
35366 övning 5
35367 övningarna 1
35368 övningsflygning 1
35369 övre 2
35370 övrig 6
35371 övriga 91
35372 övrigas 1
35373 övrigt 103
35374 – 148
