1 ! 1428
2 " 1407
3 $ 2
4 % 7
5 & 7
6 ' 21
7 ( 917
8 ) 981
9 ): 47
10 + 5
11 , 20629
12 - 1787
13 -(EN 1
14 -(ES 1
15 -54 1
16 -En 1
17 -bearbetning 1
18 -er 1
19 -företag 1
20 -kravet 1
21 -organ 3
22 -politik 1
23 -resurserna 1
24 -är 1
25 . 22976
26 .. 1
27 ... 115
28 .... 3
29 .adp 1
30 .lpk 1
31 .mdb 1
32 .odc 1
33 .udl 1
34 .xml 1
35 .xsd 1
36 .xsl-fil 2
37 / 68
38 0 1
39 0,01 3
40 0,4 1
41 0,6 1
42 0,7 4
43 00.05 1
44 000 102
45 000-3 1
46 008 2
47 0113 1
48 0550 1
49 0652 1
50 09.00 1
51 1 116
52 1,2 2
53 1,27 1
54 1,4 1
55 1,5 1
56 1,7 2
57 1,8 1
58 1,84 1
59 1,9 1
60 1-100 1
61 1-2 1
62 1-3 1
63 1-bil 1
64 1-fonderna 1
65 1-land 1
66 1-område 1
67 1-områden 1
68 1-områdena 3
69 1-området 1
70 1-region 1
71 1-regioner 2
72 1-regionerna 3
73 1-status 2
74 1-stöden 1
75 1/3 1
76 10 48
77 10,9 1
78 10.000 1
79 10.40 1
80 100 27
81 100-procentig 1
82 100c 1
83 101 1
84 101-200 1
85 102 2
86 103 2
87 104 2
88 105 4
89 106 1
90 107 3
91 107:e 1
92 108 2
93 11 33
94 11,3 1
95 11.00 11
96 11.1 3
97 11.10 1
98 11.25 1
99 11.30 7
100 110 2
101 110:e 1
102 11195/1/1999 1
103 112 1
104 11287/1/1999 1
105 112:e 1
106 114 1
107 115 1
108 116:e 1
109 119:e 1
110 11d 1
111 12 34
112 12.00 28
113 12.25 1
114 12.30 1
115 12.40 1
116 12/99 3
117 120 2
118 122 1
119 123 2
120 1244 6
121 12485/1/1999 1
122 12487/1/1999 1
123 125 1
124 1257/99 1
125 1260 1
126 1260/1999om 1
127 1260/99 1
128 127 1
129 1284 2
130 129 1
131 13 53
132 13,5 2
133 13,9 1
134 13-14 3
135 13.05 1
136 13.23 1
137 13.40 1
138 13.55 1
139 130 2
140 133.2 1
141 137 1
142 138 1
143 138.4 1
144 14 45
145 14,7 1
146 14.10 1
147 140 2
148 1408 1
149 14094/1999 2
150 142 1
151 143 1
152 1448 1
153 15 50
154 15,2 1
155 15,4 1
156 15-minuters 1
157 15.00 5
158 15.45 1
159 15.50 1
160 150 7
161 152 11
162 158 5
163 158.1 1
164 159 1
165 16 27
166 16.05 1
167 16.30 2
168 1626 1
169 1626/94 1
170 1638 1
171 164 2
172 166 2
173 167 3
174 17 18
175 17.30 1
176 170 1
177 174 1
178 1762 2
179 177 2
180 1775 1
181 178 1
182 18 29
183 18.00 4
184 180 1
185 1800-talet 2
186 1800-talets 2
187 1809 2
188 1857 1
189 1875 1
190 19 10
191 19.05 1
192 19.15 1
193 19.30 1
194 19.40 1
195 19.50 1
196 190 2
197 1900 1
198 1900-talet 4
199 1900-talets 1
200 191 1
201 1910 3
202 1917 1
203 1923 1
204 1929 3
205 193 1
206 1930-talet 2
207 194 1
208 1940 1
209 1945 1
210 1947 4
211 1948 1
212 1949 2
213 195 1
214 1952 1
215 1953 2
216 1955 1
217 1957 6
218 1958 1
219 1959 2
220 1960 2
221 1967 7
222 1969 2
223 1970 1
224 1973 4
225 1974 3
226 1975 2
227 1976 2
228 1977 2
229 1978 1
230 1979 2
231 1980-talet 2
232 1981 1
233 1982 2
234 1983 1
235 1984 4
236 1986 7
237 1987 3
238 1988 4
239 1989 6
240 1990 12
241 1990-talet 6
242 1991 5
243 1992 15
244 1993 16
245 1993-1995 2
246 1994 20
247 1994-1999 5
248 1995 24
249 1995-1997 1
250 1996 28
251 1996-1997 1
252 1997 56
253 1997/0067(COD 2
254 1997/0194(COD 2
255 1997/0352(CNS 1
256 1997/0370(COD 2
257 1997/0371(COD 2
258 1998 57
259 1998-2002 2
260 1998/0097(COD 1
261 1998/0106(COD 2
262 1998/0141 2
263 1998/0169(COD 2
264 1998/0242(COD 1
265 1998/0249(COD 1
266 1998/0324(COD 2
267 1999 154
268 1999-2000 1
269 1999-2004 1
270 1999-2006 1
271 1999/0012(COD 1
272 1999/0013(CNS 1
273 1999/0015(COD 1
274 1999/0020(COD 1
275 1999/0083 1
276 1999/0090(COD 1
277 1999/0168(CNS 2
278 1999/0196(CNS 2
279 1999/0199(CNS 2
280 1999/0218(CNS 1
281 1999/0222(CNS 1
282 1999/0224(CNS 1
283 1999/0228(CNS 1
284 1999/0240(CNS 2
285 1999/0803(CNS 1
286 1999/0805(CNS 1
287 1999/0806(CNS 1
288 1999/0809(CNS 1
289 1999/0821(CNS 2
290 1999/0825(CNS 2
291 1999/2115(COS 1
292 1999/2121(COS 2
293 1999/2123(COS 1
294 1999/2127(COS 1
295 1999/2150(COS 2
296 1999/2155(COS 2
297 1999/2182(COS 2
298 1999/2186(COS 1
299 1999/468 4
300 2 93
301 2,3 1
302 2,487 1
303 2,5 2
304 2,6 3
305 2,8 3
306 2,9 1
307 2-område 1
308 2-områdena 1
309 2-programmet 1
310 2-stöd 1
311 2.1 1
312 2.2 2
313 2.7 2
314 20 55
315 20.15 1
316 20.25 1
317 20.30 2
318 200 16
319 2000 141
320 2000- 1
321 2000-2001 1
322 2000-2004 6
323 2000-2005 8
324 2000-2006 25
325 2000-2010 1
326 2000-buggen 1
327 2000-filformat 3
328 2000-korsetten 1
329 2000-paketet 1
330 2000-platser 1
331 2000-programmet 4
332 2000-talet 5
333 2000-talets 2
334 2000-versionen 1
335 2000/2046(COS 2
336 2001 15
337 2002 35
338 2002- 2
339 2002-filformat 2
340 2003 10
341 2004 4
342 2005 4
343 2006 11
344 2007 2
345 2008 1
346 2010 10
347 2012 3
348 2020 12
349 2025 1
350 2034 1
351 205 1
352 21 16
353 21.00 5
354 21.1 1
355 21.55 1
356 2100 1
357 21:a 5
358 22 20
359 22,5 1
360 22.3 1
361 22.41 1
362 2200 1
363 226 1
364 22a 1
365 23 10
366 23,7 1
367 23-24 2
368 23.50 1
369 23.55 1
370 235- 1
371 24 21
372 24,5 1
373 240 2
374 243 1
375 245 1
376 246 1
377 248 2
378 249 4
379 25 41
380 25,7 1
381 25,9 1
382 25-åriga 1
383 250 3
384 251 1
385 255 4
386 25ºC 1
387 26 17
388 262 1
389 263 1
390 27 11
391 270 3
392 27º 1
393 28 18
394 28,2 1
395 280 4
396 280.4 1
397 28:e 1
398 29 11
399 29,9 2
400 29.4 1
401 299.2 2
402 2l:a 1
403 3 64
404 3,5 1
405 3,604 1
406 3,8 2
407 3,9 1
408 3-4 1
409 3-liter-bilar 1
410 3-liters-bilen 1
411 3.1 1
412 3.8 1
413 3/4 2
414 30 33
415 30,8 1
416 300 11
417 300.3 1
418 3062 1
419 308- 1
420 30:1 1
421 31 21
422 310 1
423 314 1
424 32 10
425 33 10
426 33,4 1
427 332 1
428 34 12
429 34.1.1 1
430 34.2 2
431 340 1
432 344 1
433 347 2
434 35 15
435 35-40 1
436 35-timmarslagen 1
437 35-timmarsvecka 1
438 35-årige 1
439 350 3
440 36 7
441 3605/93 3
442 363 2
443 366 1
444 367 1
445 37 23
446 37.2 5
447 37/60/92 1
448 370 3
449 378 2
450 38 12
451 388 2
452 39 10
453 394/2000 1
454 4 72
455 4,3 1
456 4,5 1
457 4,875 1
458 4-5 1
459 4.2 1
460 4.5 1
461 40 31
462 40-aktien 1
463 40-procentigt 1
464 400 12
465 41 8
466 410 1
467 42 8
468 42.2 1
469 42.5 1
470 43 12
471 43- 1
472 44 10
473 444 2
474 45 20
475 45-varvare 1
476 451 1
477 453 1
478 46 6
479 462 1
480 47 7
481 476 1
482 47e 1
483 48 9
484 49 8
485 4:ans 1
486 5 58
487 5,1 1
488 5,2 1
489 5,3 1
490 5,35 1
491 5,5 2
492 5,8 1
493 5-10 1
494 5.4 1
495 5.5 1
496 50 44
497 50- 1
498 50-tal 1
499 50-talskulturen 1
500 50-årsdagen 1
501 50-årsjubileum 1
502 50-årsjubiléum 1
503 500 13
504 50000 1
505 5060/1999 1
506 51 3
507 5116/1999 2
508 519 1
509 52 3
510 520 2
511 522 1
512 53 6
513 535 2
514 54 4
515 540 1
516 541 1
517 55 5
518 551 1
519 552 1
520 55:e 2
521 55º 1
522 56 5
523 56:e 3
524 57 2
525 57,5 1
526 5713/1999 1
527 58 2
528 59 4
529 5b 3
530 5b-området 1
531 6 64
532 6,07 1
533 6,4 2
534 6.1 4
535 60 21
536 60-talet 1
537 600 4
538 60:1 1
539 60º 1
540 61 1
541 613 8
542 615 1
543 62 3
544 623 2
545 63 2
546 64 1
547 65 3
548 650 1
549 6500 1
550 658 1
551 66 1
552 66,3 1
553 67 3
554 68 2
555 685/95 1
556 69 2
557 69.2 2
558 7 73
559 7,2 2
560 7,42 1
561 7,5 1
562 7-9 1
563 7.0 1
564 7.1 3
565 7.2 1
566 70 10
567 70/524 7
568 700 10
569 70:e 1
570 71 8
571 717 1
572 72 2
573 72:a 2
574 73 2
575 73,9 1
576 74 1
577 747:an 1
578 74:1 1
579 75 11
580 76 4
581 768 1
582 77 3
583 78 2
584 784 1
585 79 4
586 79/409 1
587 8 38
588 80 30
589 80-90 1
590 80-procentiga 1
591 80-talet 1
592 800 8
593 8095/1/1999 2
594 81 7
595 81(rev 1
596 81.1 5
597 81.3 5
598 82 8
599 83 3
600 830 1
601 84 2
602 85 9
603 85/611 4
604 850 9
605 850/98 1
606 86 4
607 87 5
608 87.1 1
609 87.2 1
610 88 4
611 88/591 2
612 89 3
613 9 35
614 9,2 1
615 9,5 2
616 9.00 1
617 9.1 1
618 90 17
619 90-talet 2
620 90/220 6
621 90/424 3
622 900 3
623 9085/3/1999 2
624 91 2
625 91/68 2
626 9178/1999 1
627 919 1
628 92 1
629 92/43 1
630 93 2
631 93/53 2
632 93/75 1
633 94 5
634 94/55 2
635 94/728 1
636 95 21
637 95/35 1
638 96 1
639 96/23 1
640 96/35 3
641 96/71 2
642 96/96 1
643 9614/1999 1
644 9636/1999 1
645 97 2
646 97-filformat 1
647 97/67 1
648 97/99 1
649 9767 1
650 97:e 1
651 98 3
652 99 2
653 99th 1
654 : 1053
655 ; 411
656 ? 1007
657 A 13
658 A-tjänstemän 1
659 A. 2
660 A32 1
661 A4-0029/2000 1
662 A4-0072/97 1
663 A5-0001/2000 1
664 A5-0002/2000 1
665 A5-0003/2000 2
666 A5-0004/2000 1
667 A5-0006/00 1
668 A5-0006/2000 2
669 A5-0007/2000 3
670 A5-0008/2000 3
671 A5-0009/2000 2
672 A5-0010/2000 2
673 A5-0011/2000 2
674 A5-0012/2000 2
675 A5-0013/2000 2
676 A5-0014/2000 2
677 A5-0015/2000 2
678 A5-0015/2000)av 1
679 A5-0016/2000 2
680 A5-0017/2000 3
681 A5-0018/2000 2
682 A5-0019/2000 3
683 A5-0020/2000 3
684 A5-0021/2000 2
685 A5-0022/2000 2
686 A5-0023/2000 3
687 A5-0025/2000 2
688 A5-0026/2000 1
689 A5-0027/2000 3
690 A5-0028/2000 1
691 A5-0029/2000 2
692 A5-0031/2000 3
693 A5-0032/2000 3
694 A5-0033/2000 3
695 A5-0034/2000 3
696 A5-0035/2000 1
697 A5-0036/2000 2
698 A5-0037/2000 1
699 A5-0038/2000 2
700 A5-0039/2000 1
701 A5-0040/2000 1
702 A5-0041/2000 2
703 A5-0043/2000 2
704 A5-0048/2000 1
705 A5-0051/2000 1
706 A5-0069/1999 1
707 A5-0073/1999 1
708 A5-0078/1999 1
709 A5-0087/1999 1
710 A5-0104/1999 2
711 A5-0105/1999 2
712 A5-0106/1999 1
713 A5-0107/1999 2
714 A5-0108/1999 2
715 A5­0030/2000 1
716 ABB 4
717 ABB-Alsthom 2
718 ABB-Alstom 2
719 ABC 1
720 ADOX 1
721 ADR 1
722 AKTUELLA 2
723 ALE 1
724 ALE- 1
725 ALE-gruppen 2
726 ANSI 16
727 ANSI-89 10
728 ANSI-92 11
729 ANSI-92-frågor 1
730 ANSI-92-läge 1
731 ANSI-syntax 1
732 ANVÄNDNING 1
733 ATT 1
734 AV 1
735 AVC 2
736 AVS 7
737 AVS-EU 3
738 AVS-EU-avtalet 1
739 AVS-EU-partnerskapet 1
740 AVS-EU:s 11
741 AVS-grannar 1
742 AVS-gruppen 1
743 AVS-gruppens 1
744 AVS-land 1
745 AVS-landet 1
746 AVS-länder 5
747 AVS-länderna 35
748 AVS-ländernas 9
749 AVS-partner 3
750 AVS-samarbetet 3
751 AVS-staterna 3
752 AVS-staternas 2
753 Aaron 1
754 Absaloms 1
755 Absolut 3
756 Accepterandet 1
757 Access 41
758 Access-databas 5
759 Access-databaser 2
760 Access-databasobjekt 1
761 Access-fil 2
762 Access-filen 1
763 Access-filer 1
764 Access-format 1
765 Access-projekt 4
766 Access-projektet 5
767 Act 2
768 Action 1
769 Adam 1
770 Adamson 7
771 Adana 1
772 Adapt 2
773 Adapt- 1
774 Adapt-projekt 1
775 Additionalitet 1
776 Adelaide 1
777 Adenauer 1
778 Adieu 3
779 Adjö 2
780 Administration 1
781 Administratör 1
782 Administratören 1
783 Admiral 1
784 Adolf 2
785 Adriatiska 3
786 Advanced 1
787 Adventures 1
788 Advertising 1
789 Advokaten 1
790 Afrika 53
791 Afrikanska 2
792 Afrikas 2
793 Afrodites 1
794 Agenda 21
795 Agents 1
796 Agliettas 1
797 Agrifin-rådet 1
798 Agustaaffären 1
799 Aha 1
800 Ahern 8
801 Ahmed 1
802 Ahoy 1
803 Aids 1
804 Aidsbehandlingar 1
805 Aidsproblemet 1
806 Air 2
807 Aires 1
808 Airways 1
809 Akkuyu 2
810 Akköy 1
811 Aktivera 1
812 Aktiviteterna 1
813 Alan 1
814 Alavanos 9
815 Albacète 1
816 Albaner 1
817 Albanien 13
818 Albert 1
819 Albright 1
820 Aldrig 5
821 Alex 3
822 Alexander 3
823 Alexandra 2
824 Alexandros 1
825 Alfanjurt 1
826 Alfen 1
827 Algarve 1
828 Algeriet 1
829 Algeriets 1
830 Algonquin 3
831 Alicante 2
832 Alicante-byrån 1
833 Alice 3
834 Alkartasuna 1
835 Alkoholmonopol 1
836 Alkoholpolitiken 1
837 All 4
838 Alla 88
839 Alldeles 6
840 Allen 1
841 Allesammans 1
842 Allmänheten 2
843 Allmänna 1
844 Allmänt 3
845 Allra 1
846 Allt 45
847 Alltför 3
848 Alltid 1
849 Allting 3
850 Alltsedan 3
851 Alltså 5
852 Alluvia 1
853 Almería 4
854 Alonso 1
855 Alperna 1
856 Alsace 4
857 Alsthom 1
858 Alstom 2
859 Altener 8
860 Altener-program 1
861 Altener-programmet 9
862 Alternativet 1
863 Alyssandrakis 3
864 Amadeus 1
865 Amado 4
866 Ambitionen 1
867 Ambrogio 1
868 Amerika 7
869 Amerikaner 1
870 Amerikanerna 1
871 Amerikas 5
872 Amiens 1
873 Amin 2
874 Amins 2
875 Ammokosto 1
876 Amnesty 1
877 Amoco 2
878 Amoco-Cádiz 1
879 Amoko 5
880 Amos 1
881 Amsterdam 17
882 Amsterdamfördrag 1
883 Amsterdamfördraget 46
884 Amsterdamfördragets 1
885 Amsterdamresterna 1
886 Amsterdams 1
887 Andalusien 14
888 Andelen 1
889 Andersens 1
890 Andersonbetänkandet 1
891 Andersson 19
892 Anderssonbetänkandet 3
893 Anderssons 8
894 Andliga 1
895 Andra 16
896 Andrabehandlingsrekommendation 5
897 Andrei 1
898 Andrej 14
899 Andrew 2
900 Ange 1
901 Angelilli 1
902 Angola 33
903 Angolafrågan 1
904 Angolas 2
905 Angående 57
906 Anhållandena 1
907 Ankara 5
908 Ankaras 1
909 Anledningen 2
910 Anläggning 1
911 Anmälningsplikten 1
912 Anna 2
913 Annan 1
914 Annars 10
915 Anpassa 2
916 Anpassningen 1
917 Anser 14
918 Anslagen 1
919 Anslagsbeloppet 1
920 Ansträngningarna 1
921 Anställd 1
922 Anställda 1
923 Ansvaret 4
924 Ansvarig 1
925 Ansvariga 1
926 Ansvarsfrihet 1
927 Ansvarsfriheten 1
928 Antagandet 1
929 Antal 2
930 Antalet 3
931 Antar 1
932 Antas 1
933 Antibiotika 1
934 Antingen 6
935 Antwerpen 1
936 António 3
937 Anvers 1
938 Använd 1
939 Använda 5
940 Användandet 1
941 Användare 3
942 Användaren 3
943 Användarna 2
944 Användning 1
945 Användningen 4
946 Anwar 1
947 Aparicio 1
948 Apollo 1
949 Apostrofen 1
950 Applications 1
951 Applåder 17
952 Apropå 3
953 Arabic 1
954 Arabiska 1
955 Arabrepubliken 1
956 Arabvärldens 1
957 Arafat 3
958 Arafats 2
959 Arbete 1
960 Arbetet 7
961 Arbetskultur 1
962 Arbetslöshet 1
963 Arbetslösheten 2
964 Arbetslöshetssiffrorna 1
965 Arbetsmarknad 1
966 Arbetsmarknaden 1
967 Arbetsmarknadsministeriet 1
968 Arbetspasset 1
969 Arbetsplan 2
970 Arbetsplanen 1
971 Arbetstagarna 1
972 Arbetstidsdirektivet 1
973 Arbetsvillkoren 1
974 Argumentet 1
975 Ari 1
976 Ariane 3
977 Arizona 5
978 Arkimedes 1
979 Arkiv 1
980 Arkiv-menyn 1
981 Armarna 1
982 Armenien 15
983 Arms 1
984 Arousa 1
985 Artas 1
986 Arthur 2
987 Artikel 6
988 Artikeln 1
989 Artiklarna 2
990 Arts 1
991 Asahe 4
992 Asien 4
993 Aspe-dalen 1
994 Aspects 1
995 Assad 2
996 Associations 2
997 Asturien 1
998 Ataturk-dammarna 1
999 Atatürkdammarna 1
1000 Aten 1
1001 Athen 1
1002 Athena 4
1003 Atlantalliansen 1
1004 Atlantbågens 1
1005 Atlanten 14
1006 Atlantic 1
1007 Atlantkust 1
1008 Atlantkusten 3
1009 Atlantkustens 1
1010 Att 129
1011 Attacken 1
1012 Attwool 3
1013 Attwooll 6
1014 Attwoolls 1
1015 Atxalandabaso 2
1016 Aubert 1
1017 Auerbach 2
1018 Aung 1
1019 Auroi 2
1020 Auschwitz 2
1021 Auster 35
1022 Austern 1
1023 Austers 8
1024 Australien 1
1025 Authoring 1
1026 Auto 1
1027 AutoFilter-knappen 1
1028 Autofilter 1
1029 Autofiltrering 1
1030 Auvergne 1
1031 Av 76
1032 Avbrottet 1
1033 Avbrytande 3
1034 Avenue 3
1035 Avfallet 1
1036 Avgången 1
1037 Aviano 1
1038 Avlägset 1
1039 Avreglering 2
1040 Avregleringen 2
1041 Avsaknaden 1
1042 Avsatta 1
1043 Avser 1
1044 Avsevärda 1
1045 Avsikten 3
1046 Avskaffandet 1
1047 Avslutande 1
1048 Avslutningsvis 41
1049 Avslöja 1
1050 Avtal 1
1051 Avtalen 1
1052 Avtalens 1
1053 Avtalet 9
1054 Azerbajdzjan 1
1055 Aziz 1
1056 Aznar 5
1057 Azorerna 5
1058 B 9
1059 B. 4
1060 B1-382 1
1061 B1-500 1
1062 B2-5122 1
1063 B5-0003/2000 2
1064 B5-0009/2000 2
1065 B5-0010/2000 1
1066 B5-0011/2000 1
1067 B5-0012/2000 1
1068 B5-0040/99 1
1069 B5-0041/99 1
1070 B5-0125/2000 1
1071 B5-0132/2000 1
1072 B5-0136/2000 1
1073 B5-0140/2000 1
1074 B5-0141/2000 1
1075 B5-0142/2000 1
1076 B5-0148/2000 1
1077 B5-0149/2000 1
1078 B5-0150/2000 1
1079 B5-0151/2000 1
1080 B5-0152/2000 1
1081 B5-0153/2000 1
1082 B5-0154/2000 1
1083 B5-0155/2000 1
1084 B5-0156/2000 1
1085 B5-0157/2000 1
1086 B5-0158/2000 1
1087 B5-0159/2000 1
1088 B5-0160/2000 1
1089 B5-0161/2000 1
1090 B5-0162/2000 1
1091 B5-0163/2000 1
1092 B5-0164/2000 1
1093 B5-0165/2000 1
1094 B5-0166/2000 1
1095 B5-0167/2000 1
1096 B5-0168/2000 1
1097 B5-0169/2000 1
1098 B5-0170/2000 1
1099 B5-0171/2000 1
1100 B5-0172/2000 1
1101 B5-0173/2000 1
1102 B5-0174/2000 1
1103 B5-0175/2000 1
1104 B5-0176/2000 1
1105 B5-0177/2000 1
1106 B5-0178/2000 1
1107 B5-0179/2000 1
1108 B5-0180/2000 1
1109 B5-0181/2000 2
1110 B7 1
1111 B7-0 1
1112 B7-04 1
1113 B7-4011 1
1114 B7-4012 1
1115 B7-6201 1
1116 BAT 1
1117 BBC 5
1118 BBC-intervju 1
1119 BBC:s 1
1120 BNI 13
1121 BNI-tillväxt 1
1122 BNP 9
1123 BP 1
1124 BRAY 1
1125 BRÅDSKANDE 2
1126 BSE 13
1127 BSE-epidemin 1
1128 BSE-krisen 4
1129 BSE-tester 1
1130 BSE-typ 1
1131 BSE-utskott 1
1132 BSE-utskottets 1
1133 BYRÅ 1
1134 Babitskij 15
1135 Babitskijaffären 1
1136 Babitskijs 3
1137 Baconsmörgåsarna 1
1138 Bakom 7
1139 Balfe 1
1140 Balford-förklaringen 1
1141 Balkan 51
1142 Balkanhalvöns 1
1143 Balkanländerna 2
1144 Balkanregionen 1
1145 Balkanrepublik 1
1146 Balkans 4
1147 Banantvisten 1
1148 Bandet 1
1149 Bangemann 1
1150 Bangkok 1
1151 Bank 1
1152 Bankgarantier 1
1153 Bankrutten 1
1154 Banotti 9
1155 Bara 18
1156 Barak 6
1157 Baraks 3
1158 Barcelonaprocess 1
1159 Barcelonaprocessen 1
1160 Barcelonaprocessens 1
1161 Baren 2
1162 Barents 1
1163 Baringdorf 9
1164 Barn 4
1165 Barnet 1
1166 Barnhill 1
1167 Barnier 28
1168 Barniers 4
1169 Barry 1
1170 Bartho 1
1171 Bartlebys 1
1172 Barzanti 1
1173 Barzantibetänkandet 1
1174 Barón 6
1175 Basel 1
1176 Basel-Mulhouse-flygplatsen 1
1177 Bashi 1
1178 Basic 2
1179 Basic-projektet 1
1180 Baskien 15
1181 Baskiens 2
1182 Bassam 1
1183 Basse-Normandie 1
1184 Bastille 1
1185 Battery 1
1186 Bautista 1
1187 Bay 1
1188 Bayley 6
1189 Bayley's 1
1190 Bayleys 5
1191 Bazin 1
1192 Beakta 1
1193 Beatles 3
1194 Beazley 1
1195 Bedfordshire 1
1196 Bediener 1
1197 Bedrägeri 1
1198 Bedrägeri- 1
1199 Bedömningen 2
1200 Beets 1
1201 Befolkningarnas 1
1202 Befolkningen 3
1203 Befordringssystemet 1
1204 Begreppet 2
1205 Begränsa 1
1206 Begränsningar 1
1207 Begär 1
1208 Behandlingen 2
1209 Behöver 3
1210 Bekvämlighetsflaggen 2
1211 Bekämpandet 1
1212 Bekämpning 1
1213 Belgien 16
1214 Belgiens 2
1215 Belgrad 8
1216 Belgrads 2
1217 Belize 2
1218 Belzecs 1
1219 Ben-Gurion 3
1220 Benelux 1
1221 Benenden 1
1222 Benengeli-kvartetten 1
1223 Berend 9
1224 Berendbetänkandet 1
1225 Berends 2
1226 Berenguer 3
1227 Berg 1
1228 Bergen 6
1229 Berger 11
1230 Bergerbetänkandet 1
1231 Berlin 16
1232 Berlinavtalen 1
1233 Berlinmurens 1
1234 Bern- 1
1235 Bern-konventionen 1
1236 Bernard 12
1237 Bernd 3
1238 Bernie 1
1239 Bernié 1
1240 Beroende 1
1241 Beroendet 1
1242 Beror 1
1243 Berthu 5
1244 Bertinotti 1
1245 Berätta 1
1246 Beskrivningen 1
1247 Beslut 1
1248 Besluten 1
1249 Beslutet 9
1250 Beslutsfattandet 1
1251 Besque 1
1252 Bestämmelserna 1
1253 Besättningen 1
1254 Betala 1
1255 Betoningen 1
1256 Beträffande 18
1257 Betty 1
1258 Betydande 1
1259 Betydelsen 1
1260 Betänkande 52
1261 Betänkandena 1
1262 Betänkandet 14
1263 Betänkligheterna 1
1264 Beveridges 1
1265 Beviljandet 1
1266 Beviset 2
1267 Bibel 2
1268 Bibeln 2
1269 Bidraget 1
1270 Big 5
1271 Bilbao 2
1272 Bilder 2
1273 Bilen 1
1274 Bilindustrin 1
1275 Bilkonceptet 1
1276 Bill 1
1277 Billobbyn 2
1278 Biltillverkare 2
1279 Birds 1
1280 Biscaya 1
1281 Biscayabukten 3
1282 Biscayagolfen 4
1283 Biståndet 1
1284 Biståndsgivarens 1
1285 Biståndsnivån 2
1286 Bit 1
1287 Bjerregaard 1
1288 Blak 2
1289 Blanco 3
1290 Bland 14
1291 Blanda 1
1292 Bli 1
1293 Blok 1
1294 Blokland 1
1295 Blooms 1
1296 Blotts 1
1297 Blums 1
1298 Blåfenad 1
1299 Boetticher 1
1300 Bohéme 1
1301 Boken 1
1302 Bokhållaren 1
1303 Bokläsare 1
1304 Bolaget 2
1305 Bolagets 2
1306 Bolagsdirektören 1
1307 Bolkestein 19
1308 Bolkesteins 1
1309 Bologna 1
1310 Bom 1
1311 Bomber 1
1312 Bonde 7
1313 Bonino 2
1314 Bonino-listan 1
1315 Booz 1
1316 Bor 1
1317 Borde 8
1318 Bordeaux 1
1319 Borgia 1
1320 Borgin 6
1321 Borgins 2
1322 Borràs 3
1323 Bortanför 1
1324 Bortom 4
1325 Bortre 1
1326 Bortsållning 1
1327 Bos 1
1328 Bosnien 5
1329 Bosnien-Hercegovina 1
1330 Bosnien-Herzegovina 4
1331 Bosniens 1
1332 Bosse 1
1333 Boston 1
1334 Bosättarna 1
1335 Botswana 1
1336 Bourlanges 6
1337 Bouwman 10
1338 Bowe 2
1339 Bowis 2
1340 Boyne 3
1341 Boynes 2
1342 Boynesmynningen 1
1343 Boynesmynningens 1
1344 Bra 3
1345 Braer 2
1346 Braerkatastrofen 1
1347 Brahim 1
1348 Brandenburg 2
1349 Branschen 1
1350 Brasilien 3
1351 Bravery 1
1352 Bray 41
1353 Bredden 1
1354 Bremen 1
1355 Brempt 1
1356 Bresjnevs 1
1357 Bretagne 16
1358 Bretagnes 3
1359 Bretonne 1
1360 Brevbäraren 1
1361 Brevet 1
1362 Brian 1
1363 Brist 2
1364 Bristen 1
1365 Bristerna 1
1366 British 3
1367 Brittan 1
1368 Brittiska 1
1369 Broadway 4
1370 Broek 1
1371 Brok 18
1372 Brokbetänkandet 2
1373 Broks 4
1374 Bronislav 1
1375 Brottsligheten 1
1376 Brovina 8
1377 Brovinas 1
1378 Brown 1
1379 Brundtland-rapporten 1
1380 Bruno 1
1381 Bryssel 54
1382 Bryssel-I 1
1383 Bryssel-II 1
1384 Brysselartikeln 1
1385 Brysselbyråkrater 1
1386 Brysselbyråkratin 1
1387 Brysselfederalistiskt 1
1388 Brysselfördraget 1
1389 Bryssels 2
1390 Brysselteknokraternas 1
1391 Bränningens 1
1392 Bröderna 1
1393 Budapest 3
1394 Budget- 1
1395 Budgetförordningen 2
1396 Budgetmedlen 1
1397 Budgetplanerna 1
1398 Budgetutskottet 1
1399 Buenos 1
1400 Buesa 5
1401 Building 1
1402 Bulgarien 8
1403 Bull 1
1404 Bundestag 1
1405 Burkes 2
1406 Burkina 1
1407 Burma 11
1408 Burrow 2
1409 Bush 1
1410 Busquin 1
1411 Busquins 2
1412 Bygget 1
1413 Byn 1
1414 Byrne 11
1415 Byrån 7
1416 BÄTTRE 1
1417 Bägge 1
1418 Bär 1
1419 Bästa 1
1420 Bäste 2
1421 Bättre 1
1422 Båda 10
1423 Både 8
1424 Béguin 2
1425 Böcker 1
1426 Böge 6
1427 Böges 2
1428 Böhm 1
1429 Bör 1
1430 Börja 1
1431 Bösch 1
1432 Bülent 2
1433 C 5
1434 C. 4
1435 C4-0018/98 1
1436 C4-0026/1999 2
1437 C4-0212/1999 1
1438 C4-0350/1998 1
1439 C4-0351/1998 1
1440 C4-0352/1999 1
1441 C4-0465/1998 1
1442 C4-0497/98-98/0126 1
1443 C4-0715/98-98/0318(SYN 1
1444 C5-0004/1999 1
1445 C5-0013/2000 1
1446 C5-0014/00 1
1447 C5-0020/1999 1
1448 C5-0040/2000 1
1449 C5-0045/00 1
1450 C5-0045/2000 1
1451 C5-0050/2000 1
1452 C5-0069/1999 1
1453 C5-0081/2000 2
1454 C5-0091/1999 1
1455 C5-0095/1999 1
1456 C5-0112/1999 1
1457 C5-0120/99 1
1458 C5-0122/1999 1
1459 C5-0134/1999 2
1460 C5-0156/1999 2
1461 C5-0166/1999 2
1462 C5-0167/1999 1
1463 C5-0174/1999 2
1464 C5-0176/1999 2
1465 C5-0180/1999 2
1466 C5-0208/1999 2
1467 C5-0209/1999 2
1468 C5-0222/1999 2
1469 C5-0251/99 1
1470 C5-0253/1999 2
1471 C5-0260/1999 1
1472 C5-0302/1999 1
1473 C5-0303/1999 1
1474 C5-0305/1999 1
1475 C5-0308/1999 2
1476 C5-0323/99 1
1477 C5-0327/1999 2
1478 C5-0331/1999 1
1479 C5-0332/1999 2
1480 C5-0333/1999 2
1481 C5-0334/1999 2
1482 C5-0341/1999 2
1483 CAC 3
1484 CECAF:s 1
1485 CEN 8
1486 CEN:s 4
1487 CERN 1
1488 CIA 3
1489 CIP 1
1490 CNS 1
1491 COD 1
1492 COPA 1
1493 CORUS 1
1494 COSV 1
1495 CSS 3
1496 CSS-fil 2
1497 CSU-gruppens 1
1498 CSU:s 2
1499 CTRL-C. 1
1500 CTRL-V. 1
1501 Cabrols 1
1502 Cadiz 4
1503 Cadiz-katastrofen 2
1504 Cadou 1
1505 Caesarea 1
1506 Caillaux 1
1507 Calais 1
1508 Cambridge 1
1509 Camdessus 1
1510 Campos 1
1511 Camre 1
1512 Camus 1
1513 Canada 1
1514 Candutyp 1
1515 Canyon 3
1516 Canyons 1
1517 Cappuccino 1
1518 Capra 1
1519 Cara-programmet 1
1520 Cardiff 2
1521 Cardiffprocessen 2
1522 Carlo 1
1523 Caroline 1
1524 Casablanca 1
1525 Casaca 1
1526 Casas 2
1527 Cascading 1
1528 Cashman 1
1529 Castro-regimen 1
1530 Caudron 1
1531 Cavalese 1
1532 Cederschiöld 13
1533 Cederschiöldbetänkandet 1
1534 Cederschiölds 5
1535 Celsius 3
1536 Cem 1
1537 Central 1
1538 Central- 11
1539 Centralamerika 2
1540 Centralasiatiska 2
1541 Centralasien 3
1542 Centralasiens 1
1543 Centralbanken 3
1544 Centralbankschefen 1
1545 Centraleuropa 2
1546 Cermis 1
1547 Cervantes 1
1548 Ceyhun 1
1549 Champagne-Ardennes 1
1550 Chanel 1
1551 Change 1
1552 Chapmanfyren 1
1553 Charente 1
1554 Charles 1
1555 Charlie 2
1556 Charlotte 1
1557 Charm 1
1558 Chefen 1
1559 Chevènement 1
1560 Chicago 3
1561 Chief 1
1562 Chile 2
1563 Chiquita 1
1564 Chissano 1
1565 Chris 1
1566 Christine 1
1567 Christopher 4
1568 Church 1
1569 Ciampi-gruppen 1
1570 Circa 1
1571 Cirka 2
1572 Cisterna 6
1573 Cisternen 1
1574 Clare 1
1575 Claude 3
1576 Clintons 1
1577 Clough 1
1578 Clément 1
1579 Coca 1
1580 Cocilovo 1
1581 Coco 1
1582 Cocoon 1
1583 Coelho 1
1584 Coffee 1
1585 Cohn-Bendit 6
1586 Cola 1
1587 Colombia 2
1588 Colonial 1
1589 Comartkommitté 1
1590 Comartkommittén 1
1591 Comet 1
1592 Comité 1
1593 Commission 2
1594 Community 1
1595 Company 1
1596 Companys 1
1597 Compensation 1
1598 Components 5
1599 Components-element 1
1600 Compostela 1
1601 Compson 1
1602 Compsons 1
1603 Conakry 1
1604 Confederation 1
1605 Connaught 1
1606 Connection 1
1607 ConnectionFile 4
1608 ConnectionString 6
1609 Consortium 3
1610 Constabulary 1
1611 Contre 1
1612 Copeland 3
1613 Copyright 1
1614 Corbett 7
1615 Core-projektet 1
1616 Corinne 1
1617 Cork 3
1618 Cornelissen 1
1619 Cornwall 1
1620 Corporate 1
1621 Corpus 1
1622 Corrie 17
1623 Corrie-betänkandet 1
1624 Corriebetänkandet 1
1625 Corriebetänkandets 1
1626 Cossutta 1
1627 Costa 11
1628 Council 1
1629 Coupe 1
1630 Cox 9
1631 Coûteaux 1
1632 Crab 1
1633 Crespo 2
1634 Crespos 2
1635 Cresson 2
1636 Crisex 1
1637 Crowley 3
1638 Cummings 3
1639 Cunard 2
1640 Cunardbolaget 1
1641 Cunards 1
1642 Cunha 1
1643 Cunhabetänkandet 1
1644 Cunhas 1
1645 Curie-stipendier 1
1646 Curtis 3
1647 Curveting 1
1648 Cushnahan 1
1649 Cusí 1
1650 Cusís 2
1651 Cuxhaven 1
1652 Cyaniden 1
1653 Cymru 1
1654 Cypern 74
1655 Cypernfrågan 6
1656 Cypernkonflikten 1
1657 Cypernproblemet 1
1658 Cyperns 14
1659 Cypernsamtalen 1
1660 Cyprian 2
1661 D 2
1662 DA 12
1663 DB-datakälla 1
1664 DB-datakällor 1
1665 DDR 1
1666 DE 14
1667 DEAF 1
1668 DEBATT 2
1669 DINA 1
1670 DISTINCT 1
1671 Da 3
1672 Dagen 1
1673 Dagens 8
1674 Dagerns 1
1675 Dagligen 3
1676 Dagmar 1
1677 Dagordningen 1
1678 Daily 1
1679 Daladiers 1
1680 Dalai 7
1681 Dalmau 1
1682 Dam 3
1683 Damaskus 3
1684 Damer 1
1685 Dando 25
1686 Dandos 3
1687 Dandy-Roly 1
1688 Daniel 8
1689 Danmark 44
1690 Danmarks 2
1691 Danny 1
1692 Dansarna 1
1693 Dansetteskivspelare 1
1694 Darmstadt 1
1695 Data 3
1696 Datablad 1
1697 Databladsläge 1
1698 Datum 1
1699 Datum- 1
1700 David 11
1701 Davids 1
1702 Davies 4
1703 Davis 2
1704 Dayton 2
1705 De 540
1706 Dead 1
1707 Debatten 5
1708 Debatterna 1
1709 Decourrière 7
1710 Decourrièrebetänkandet 1
1711 Decourrières 3
1712 Decree 1
1713 Definitionerna 1
1714 Definitivt 1
1715 Deklarationen 1
1716 Delat 1
1717 Delegationerna 1
1718 Dell'Alba 1
1719 Delningen 1
1720 Delors 8
1721 Delorskommissionens 1
1722 Delorsplanen 1
1723 Dels 2
1724 Deltagandet 1
1725 Delvis 2
1726 Dem 1
1727 Deminimus-bestämmelserna 1
1728 Demokrati 1
1729 Demokratiska 1
1730 Demonstranterna 1
1731 Den 655
1732 Denktash 2
1733 Denna 149
1734 Denne 2
1735 Deptford 1
1736 Deras 14
1737 Derbyshire 1
1738 Derivatmarknaden 1
1739 Derrick 1
1740 Desama 2
1741 Design-vyn 2
1742 Desktop 2
1743 Dess 7
1744 Dessa 126
1745 Dessert 1
1746 Dessutom 96
1747 Destabiliseringen 1
1748 Desto 3
1749 Det 2842
1750 Detaljerad 1
1751 Detaljerna 1
1752 Detaljområde 1
1753 Detektivbyrå 1
1754 Detsamma 3
1755 Detta 594
1756 Deutsche 3
1757 Developer 1
1758 Devon 1
1759 Di 14
1760 Diagongränden 2
1761 Diagram 2
1762 Dialog 2
1763 Diamantopoulou 7
1764 Dick 1
1765 Dig 1
1766 Digital 1
1767 Dimitrakopoulos 5
1768 Din 1
1769 Dineh 7
1770 Dinehbefolkningen 1
1771 Dinehindianerna 1
1772 Dinky-leksaker 1
1773 Dior 1
1774 Dipecho 1
1775 Dipechos 2
1776 Diplomatiska 1
1777 Direktivet 18
1778 Direktivets 2
1779 Direktören 1
1780 Diskrimineringen 1
1781 Diskussionen 3
1782 Diskussionens 1
1783 Diskussionsämnet 1
1784 Diskuteras 1
1785 Dit 2
1786 Dixon 1
1787 Djupare 1
1788 Dobby 12
1789 Dobbys 1
1790 Dock 13
1791 Dokumenten 1
1792 Dokumentet 2
1793 Dolorosa 1
1794 Dom 4
1795 Domarna 1
1796 Dominique 3
1797 Domstolen 2
1798 Domstolens 2
1799 Don 9
1800 Donau 17
1801 Donaus 4
1802 Donnay 1
1803 Doris 2
1804 Dorothy 1
1805 Dos 3
1806 Dostoevski 2
1807 Dostoevski's 1
1808 Doyles 1
1809 Doñana 2
1810 Doñana-katastrofen 1
1811 Dra 1
1812 Draco 8
1813 Drake 1
1814 Dreyfus-affärens 1
1815 Dricka 1
1816 Drive 7
1817 Drogheda 5
1818 Drug 1
1819 Dröjsmålet 1
1820 Drömmen 1
1821 Du 84
1822 Dubbelt 1
1823 Dublin 5
1824 Dublinfonden 1
1825 Dublinkonventionen 2
1826 Dublinkonventionerna 1
1827 Duc 1
1828 Dudley 19
1829 Dudleys 2
1830 Duhamels 1
1831 Duisenberg 3
1832 Duktig 1
1833 Dumbledore 1
1834 Dumpning 2
1835 Dunn 1
1836 Dupuis 4
1837 Dur 1
1838 Durban 1
1839 Dursley 9
1840 Dursleys 17
1841 Dutroux 1
1842 Dutroux-affären 1
1843 Dvs. 2
1844 Där 49
1845 Därav 4
1846 Därefter 14
1847 Däremot 26
1848 Därför 302
1849 Däri 1
1850 Därifrån 1
1851 Därigenom 5
1852 Därmed 17
1853 Därtill 1
1854 Därute 1
1855 Därutöver 2
1856 Därvid 3
1857 Då 65
1858 Démocratique 1
1859 Díez 5
1860 Död 1
1861 Döda 2
1862 Dörrarna 1
1863 Dührkop 3
1864 E-kolibakteriesmittat 1
1865 ECB 2
1866 ECHO 13
1867 ECHO:s 1
1868 ECHR 2
1869 ECTAA 1
1870 EDD 3
1871 EDD-Gruppen 1
1872 EDD-gruppens 3
1873 EDF-medlens 1
1874 EDU:s 1
1875 EE 2
1876 EEC 1
1877 EEG 12
1878 EFTA:s 1
1879 EG 26
1880 EG-Israel 3
1881 EG-biståndet 1
1882 EG-direktiv 2
1883 EG-direktiven 2
1884 EG-direktivet 1
1885 EG-domstolen 25
1886 EG-domstolens 3
1887 EG-fördraget 9
1888 EG-kort 9
1889 EG-kortet 7
1890 EG-obligationer 1
1891 EG-rätt 2
1892 EG-rätten 1
1893 EG-verksamheter 1
1894 EG:s 8
1895 EIF 2
1896 EKSG 2
1897 EKSG-fördraget 6
1898 EL 9
1899 ELDR 3
1900 ELDR-gruppen 3
1901 ELDR:s 1
1902 EMU 3
1903 EMU-anpassningens 1
1904 EMU-anslutning 1
1905 EMU-eran 1
1906 EMU-fördraget 1
1907 EMU-kriterierna 2
1908 EMU-medlemsstater 1
1909 EMU-projekt 1
1910 EMU-projektet 1
1911 EMU-projektets 1
1912 EMU-samarbetet 1
1913 EMU:s 5
1914 EN 75
1915 ENS 10
1916 EPP-DE 1
1917 ERUF 1
1918 ES 7
1919 ETA 8
1920 ETA-förhandlare 1
1921 ETA:s 2
1922 EU 217
1923 EU- 2
1924 EU-AVS-avtalet 1
1925 EU-AVS-sammanhanget 1
1926 EU-Medelhavsområdet 1
1927 EU-anslutningen 1
1928 EU-behörighet 1
1929 EU-beslut 1
1930 EU-bistånd 1
1931 EU-biståndet 1
1932 EU-budgeten 1
1933 EU-enheten 1
1934 EU-fonder 1
1935 EU-fördrag 2
1936 EU-fördragen 1
1937 EU-fördraget 8
1938 EU-företag 2
1939 EU-förordningar 1
1940 EU-genomsnittet 1
1941 EU-initiativ 1
1942 EU-insatser 1
1943 EU-institutioner 1
1944 EU-institutionerna 4
1945 EU-institutionernas 2
1946 EU-kandidater 1
1947 EU-kommissionen 2
1948 EU-kort 2
1949 EU-kortet 2
1950 EU-kriterierna 1
1951 EU-lagstiftningen 4
1952 EU-landet 1
1953 EU-länder 7
1954 EU-länderna 6
1955 EU-ländernas 1
1956 EU-mantra 1
1957 EU-marknaden 1
1958 EU-marknader 1
1959 EU-medborgare 5
1960 EU-medborgarnas 1
1961 EU-medel 2
1962 EU-medlemmar 2
1963 EU-medlemmarna 2
1964 EU-medlemskap 2
1965 EU-medlemsstaterna 3
1966 EU-medlemsstaternas 1
1967 EU-miljöreglerna 1
1968 EU-nivå 6
1969 EU-nivån 1
1970 EU-omfattande 1
1971 EU-ordförandeskapets 1
1972 EU-organ 2
1973 EU-pass 3
1974 EU-perspektiv 1
1975 EU-politik 1
1976 EU-program 2
1977 EU-regeringar 1
1978 EU-regi 1
1979 EU-reglerad 1
1980 EU-resurser 1
1981 EU-räntor 1
1982 EU-rätt 1
1983 EU-rättskipning 1
1984 EU-rådets 1
1985 EU-samarbetet 1
1986 EU-skeptiker 1
1987 EU-staterna 1
1988 EU-staternas 1
1989 EU-straffrätt 1
1990 EU-strukturfonder 1
1991 EU-system 1
1992 EU-sändebud 2
1993 EU-texterna 1
1994 EU-utvidgning 1
1995 EU-världen 1
1996 EU:s 125
1997 EUF 8
1998 EUF-medel 1
1999 EUF-medlen 1
2000 EUGFJ 4
2001 EUGFJ:s 1
2002 East 1
2003 Ecemis-förkastningslinjen 1
2004 Ecevit 2
2005 Echelon 3
2006 Echelon-nätet 1
2007 Edinburgh 3
2008 Editor 1
2009 Edouard 2
2010 Edward 4
2011 Edwards 4
2012 Effekten 3
2013 Effekterna 1
2014 Effektiv 2
2015 Effektiva 1
2016 Effektivitet 1
2017 Effektiviteten 2
2018 Eftarløn 2
2019 Efter 55
2020 Efterskalven 1
2021 Eftersom 75
2022 Efteråt 3
2023 Egeiska 1
2024 Egenskaper 1
2025 Egentligen 7
2026 Egypten 5
2027 Ehud 2
2028 Eichelberger 4
2029 Eichelbergers 1
2030 Eieck 1
2031 Einstein 1
2032 Ejido 26
2033 Ejidos 2
2034 Ekofin 2
2035 Ekofin-ministrar 1
2036 Ekofin-ministrarna 1
2037 Ekofin-rådet 8
2038 Ekologiskt 1
2039 Ekonomer 1
2040 Ekonomierna 1
2041 Ekonomin 4
2042 Ekonomisk 1
2043 Ekonomiska 6
2044 Ekonomistyrningen 1
2045 El 28
2046 Elbe 1
2047 Elden 1
2048 Elektriskt 1
2049 Elementen 1
2050 Elf 1
2051 Elfenbenskusten 1
2052 Elie 1
2053 Eline 1
2054 Elisabeth 1
2055 Eller 17
2056 Elles 3
2057 Elly 1
2058 Elmar 4
2059 Elorza 2
2060 Elst 1
2061 Elva 1
2062 Emellanåt 1
2063 Emellertid 12
2064 Emergency 1
2065 Emilia-Romagna 1
2066 Empire 1
2067 Employment 1
2068 Employment-initiativen 1
2069 Emprego 1
2070 Empress 1
2071 En 308
2072 Enbart 2
2073 End 1
2074 Enda 1
2075 Endast 20
2076 Eneko 1
2077 Energisituationen 1
2078 Enfopol 1
2079 Engagemang 1
2080 Engelska 2
2081 Engelsmän 1
2082 Engine 2
2083 England 11
2084 Englands 1
2085 Enigheten 1
2086 Enkelt 1
2087 Enligt 81
2088 Enorma 1
2089 Enrique 3
2090 Entebbe 1
2091 Enterprise 1
2092 Entitet 1
2093 Equal 24
2094 Equal- 1
2095 Equal-betänkande 1
2096 Equal-betänkandet 10
2097 Equal-initiativet 19
2098 Equal-initiativets 2
2099 Equal-programmet 6
2100 Equal-programmets 1
2101 Equqal 2
2102 Er 8
2103 Era 4
2104 Erebus 1
2105 Erfarenheten 4
2106 Erfarenheter 1
2107 Erfarenheterna 4
2108 Ericsson 1
2109 Erika 44
2110 Erika-katastrofen 3
2111 Erika-katastrofer 1
2112 Erika-olyckan 1
2113 Erikas 14
2114 Erith 1
2115 Eritrea 1
2116 Erkki 2
2117 Ermua 1
2118 Eros 1
2119 Errols 1
2120 Ert 7
2121 Escola 1
2122 Essen 1
2123 Essex 1
2124 Essex-Suffolk-Norfolkkusten 1
2125 Essexmaderna 1
2126 Estland 1
2127 Etiopien 6
2128 Etnisk 1
2129 Ett 152
2130 Etthundratjugotvå 1
2131 Eugene 1
2132 Euratom 4
2133 Euratomfördraget 1
2134 Euro 1
2135 Euro-Atlantiska 1
2136 Euro-Paper 1
2137 Euro-rådet 1
2138 Eurodac 4
2139 Eurodac-systemet 1
2140 Eurojust 6
2141 Euroland 3
2142 Euron 2
2143 Eurons 3
2144 Europa 711
2145 Europa-Afrika 1
2146 Europa-Medelhavsländerna 1
2147 Europademokrater 14
2148 Europademokraterna 2
2149 Europademokraternas 1
2150 Europadomstolen 1
2151 Europafrågan 1
2152 Europafrågor 1
2153 Europagrupp 1
2154 Europakonventionen 2
2155 Europaminister 2
2156 Europaministerns 1
2157 Europanivå 1
2158 Europaparlament 3
2159 Europaparlamentarikerna 1
2160 Europaparlamentet 290
2161 Europaparlamentets 118
2162 Europaparlamentsledamöternas 2
2163 Europarådet 2
2164 Europas 131
2165 Europaskatt 1
2166 Europatrupp 1
2167 Europaval 3
2168 Europavalen 4
2169 Europavalet 1
2170 Europavänligt 1
2171 Europe 4
2172 European 2
2173 Europeisk 1
2174 Europeiska 1197
2175 Europol 18
2176 Europolavtalet 1
2177 Europolkonventionen 1
2178 Europols 4
2179 Européerna 1
2180 Euroskeptikerna 1
2181 Eurostat 3
2182 Euskal 2
2183 Eusko 1
2184 Evans 7
2185 Evelyn 5
2186 Evelyns 1
2187 Eventuellt 2
2188 Exakt 1
2189 Excel 13
2190 Exceptionellt 1
2191 Exempel 6
2192 Exempelvis 2
2193 Exemplen 1
2194 Exemplet 2
2195 Experimental 1
2196 Experterna 3
2197 Expertutfrågningarna 1
2198 Explorer 3
2199 Exportera 6
2200 Expresso 1
2201 Extensible 3
2202 Exxon 3
2203 F 1
2204 F. 1
2205 FBI 2
2206 FEO 3
2207 FFP 1
2208 FFP:s 1
2209 FI 1
2210 FIPOL 1
2211 FMI 1
2212 FN 17
2213 FN-embargot 1
2214 FN-finansieringen 1
2215 FN-flyktingar 1
2216 FN-länder 1
2217 FN-närvaro 1
2218 FN-programmet 1
2219 FN-stadgan 1
2220 FN-stöd 1
2221 FN-uppdragets 1
2222 FN:s 36
2223 FPÖ 13
2224 FPÖ-ledaren 1
2225 FPÖ-medlemmar 1
2226 FPÖ:s 4
2227 FR 57
2228 FROM 1
2229 FRÅGOR 2
2230 FTSE 1
2231 FUF 1
2232 FYROM 8
2233 FYROM:s 4
2234 Fackföreningarna 1
2235 Fackföreningsrepresentanter 2
2236 Factortame-fallet 1
2237 Faim 1
2238 Fakta 2
2239 Faktum 12
2240 Fallet 5
2241 Falska 1
2242 Falskmyntning 1
2243 Falskt 1
2244 Falun 1
2245 Familjejordbruket 1
2246 Fan 1
2247 Fanns 1
2248 Far 10
2249 Farbror 2
2250 Farligt 1
2251 Farmor 5
2252 Farouk 1
2253 Fartyget 4
2254 Fartygets 1
2255 Fartygsbränslet 1
2256 Fascismen 1
2257 Faslane 2
2258 Faso 1
2259 Fast 7
2260 Fastän 1
2261 Fattas 1
2262 Fattigbasaren 1
2263 Fattigdomen 1
2264 Fattigdomsbekämpning 1
2265 Faulkner 2
2266 Fay 1
2267 Federal 1
2268 Federation 1
2269 Feira 3
2270 Felaktigt 1
2271 Felet 1
2272 Fem 6
2273 Femte 1
2274 Femton 1
2275 Femårsprogrammet 1
2276 Ferber 1
2277 Fernando 5
2278 Fernández 4
2279 Ferte 1
2280 Festmåltider 1
2281 Festus 3
2282 Festus' 1
2283 Fidji-öarna 1
2284 Field 1
2285 Filen 1
2286 Filter 1
2287 Filterfält 1
2288 Filterinställningar 1
2289 Filtrera 4
2290 Filtrerad 1
2291 Filtrerat 1
2292 Filtreringseffekter 1
2293 Filtreringsmetoder 1
2294 Fina 1
2295 Finansiella 1
2296 Finansiellt 1
2297 Finansiering 1
2298 Finansieringen 3
2299 Finansministrarna 1
2300 Fingrarna 1
2301 Finisterre 1
2302 Finland 27
2303 Finlands 1
2304 Finnarna 1
2305 Finner 2
2306 Finns 28
2307 Firman 1
2308 Fischler 18
2309 Fischlers 3
2310 Fishing 1
2311 Fisk 1
2312 Fiskare 1
2313 Fiskarnas 1
2314 Fiske 1
2315 Fiskeflottan 1
2316 Fiskeriförvaltning 3
2317 Fiskeriindustrin 1
2318 Fiskerisektorerna 1
2319 Fisket 2
2320 Fitousi 1
2321 Fitzsimons 1
2322 Fjolårets 1
2323 Fjorton 1
2324 Fjortonåriga 1
2325 Flandern 4
2326 Flats 1
2327 Flautre 1
2328 Flautres 1
2329 Fleet 1
2330 Fleetwood 1
2331 Fler 2
2332 Flera 11
2333 Flertalet 1
2334 Flexibilitet 1
2335 Flickan 3
2336 Floden 2
2337 Floderna 1
2338 Flora 8
2339 Floras 1
2340 Florenz 19
2341 Florenzbetänkandet 1
2342 Flourish 1
2343 Flugorna 1
2344 Flyg 1
2345 Flyg- 1
2346 Flygvärdinnorna 1
2347 Flytta 4
2348 Flyttfåglar 1
2349 Flämtande 1
2350 Flåsande 1
2351 Fléchard-affären 1
2352 FoU 1
2353 FoU-ramprogrammet 1
2354 Fodertillsatser 1
2355 Fog 1
2356 Folk 6
2357 Folkets 2
2358 Folkfronten 1
2359 Folkmordet 1
2360 Folkrepubliken 2
2361 Folkvalda 1
2362 Fondföretag 2
2363 Fondföretagen 1
2364 Fondsparande 1
2365 Fontaine 7
2366 Fontaines 1
2367 Food 1
2368 Force 1
2369 Ford 1
2370 Forest 1
2371 Forestier 1
2372 Formulär 1
2373 Forskarna 1
2374 Forskningen 1
2375 Forsyth 1
2376 Forsyth-Byggen 1
2377 Fort 1
2378 Fortfarande 2
2379 Fortsätt 1
2380 Fortunas 1
2381 Fotografier 1
2382 Fraga 1
2383 Fraisse 1
2384 Fram 4
2385 Framför 11
2386 Framförallt 2
2387 Framgångarna 1
2388 Framläggandet 1
2389 Framsteg 1
2390 Framstegen 2
2391 Framställningar 1
2392 Framtagandet 1
2393 Framtida 1
2394 Framtiden 1
2395 Framåt 1
2396 France 2
2397 Frances 1
2398 Francis 3
2399 Franco 2
2400 Franklin 1
2401 Frankrike 64
2402 Frankrikes 10
2403 Franoise 1
2404 Fransmännen 3
2405 Franz 3
2406 François 1
2407 Frassoni 11
2408 Fred 21
2409 Freden 1
2410 Frederiksen 1
2411 Freds 1
2412 Freds- 2
2413 Fredsprocessen 4
2414 Free 1
2415 Freetown 1
2416 Freud 1
2417 Fricks 1
2418 Frid 1
2419 Frihet 3
2420 Friheten 1
2421 Frihetspartiet 3
2422 Frihetspartiets 1
2423 Fritt 1
2424 FrontPage 2
2425 Frontera 1
2426 Fru 214
2427 Fruteau 3
2428 Främjande 2
2429 Främjandet 1
2430 Främst 2
2431 Fråga 51
2432 Frågan 46
2433 Frågestund 4
2434 Frågor 6
2435 Frågorna 5
2436 Från 21
2437 Frånvaron 1
2438 Fukuyama 1
2439 Full 2
2440 Fund 4
2441 Fundera 1
2442 Fungerar 1
2443 Funktionen 1
2444 Fy 1
2445 Fyra 4
2446 Fyrtio 1
2447 Fysiska 1
2448 Fältpil 1
2449 Fältpilen 1
2450 Färden 1
2451 Färg 1
2452 Färre 1
2453 Fästning 1
2454 Få 2
2455 Fågeln 1
2456 Får 16
2457 Följaktligen 8
2458 Följande 4
2459 Följden 3
2460 Följderna 2
2461 För 591
2462 Förbaskade 1
2463 Förbaskat 1
2464 Förbereda 1
2465 Förberedelserna 1
2466 Förbindelserna 1
2467 Förbrukningen 1
2468 Förbud 2
2469 Förbundskansler 1
2470 Förbundsrepubliken 5
2471 Fördelar 1
2472 Fördelarna 1
2473 Fördelen 2
2474 Fördomar 1
2475 Fördragen 2
2476 Fördraget 9
2477 Fördragets 1
2478 Före 8
2479 Förebyggande 2
2480 Föredragande 2
2481 Föredraganden 15
2482 Föredragandens 3
2483 Föredragningslista 3
2484 Föregående 1
2485 Förekommer 1
2486 Föreliggande 1
2487 Förenade 44
2488 Förenligheten 1
2489 Förenta 118
2490 Föresatsen 1
2491 Föreslagna 1
2492 Föreslå 1
2493 Föreställer 1
2494 Föreställningen 1
2495 Företag 2
2496 Företrädaren 1
2497 Företrädarna 1
2498 Förfalskningar 1
2499 Förfarande 1
2500 Förfarandena 1
2501 Förfarandet 3
2502 Förflyttningen 1
2503 Förhandlingar 1
2504 Förhandlingen 1
2505 Förhindra 1
2506 Förhoppningar 1
2507 Förhoppningarna 2
2508 Förhoppningen 1
2509 Förhoppningsvis 4
2510 Förintelsekonferensen 1
2511 Förintelsen 2
2512 Förklaringen 1
2513 Förlisningen 1
2514 Förlorare 1
2515 Förlusterna 1
2516 Förlåt 2
2517 Förmodligen 3
2518 Förnyelsen 1
2519 Förordningen 4
2520 Förordningens 2
2521 Förorenaren 2
2522 Förpackningar 1
2523 Förr 1
2524 Förra 8
2525 Förresten 1
2526 Församlingarna 1
2527 Försiktighet 1
2528 Försiktighetsprincipen 2
2529 Förskjutningen 1
2530 Förslag 5
2531 Förslagen 5
2532 Förslaget 14
2533 Förslagets 1
2534 Förslagsrätt 1
2535 Först 61
2536 Första 3
2537 Förstainstansrätten 1
2538 Förstelning 1
2539 Förstå 1
2540 Förståeligt 1
2541 Förstår 3
2542 Förstörelsen 1
2543 Försvarsmakten 1
2544 Försämrar 1
2545 Försåvitt 1
2546 Försök 1
2547 Försöken 1
2548 Försöket 1
2549 Förtalet 1
2550 Förteckningen 2
2551 Förtjänster 1
2552 Förtroendet 1
2553 Förtrollad 1
2554 Förutom 13
2555 Förutsatt 2
2556 Förvaltningen 2
2557 Förvaltningsbolag 1
2558 Förvisso 5
2559 Förväntningarna 1
2560 Förvärrad 1
2561 Förändring 1
2562 Förändringar 3
2563 Förändringarna 2
2564 G8-mötet 1
2565 GA-stöd 1
2566 GAL 2
2567 GASP 1
2568 GATS-avtalen 1
2569 GATT 1
2570 GATT-avtalet 2
2571 GATT-förhandlingarna 1
2572 GATT:s 1
2573 GD 1
2574 GFP 1
2575 GJP 4
2576 GJP-reformerna 1
2577 GMO 16
2578 GMO-fri 1
2579 GRANT 1
2580 GUE 3
2581 GUSP 6
2582 GYLLENROY 1
2583 Gaeta 1
2584 Gai-Hinnom 4
2585 Gala 2
2586 Galaprovinsen 1
2587 Galas 1
2588 Galeote 4
2589 Galicien 6
2590 Gallagher 4
2591 Gallaghers 2
2592 Gallierna 1
2593 Gama 3
2594 Gamla 1
2595 Gammal 1
2596 Ganska 1
2597 Garanterandet 1
2598 García 1
2599 García-Margallo 2
2600 Garcías 1
2601 Gargani 5
2602 Gascognebukten 1
2603 Gasòliba 1
2604 Gatornas 1
2605 Gaulles 1
2606 Gaza 5
2607 Gazaregionen 1
2608 Gazaremsan 2
2609 Ge 3
2610 Gehenna 1
2611 Gemelli 1
2612 Gemensam 3
2613 Gemensamma 1
2614 Gemensamt 7
2615 Gemenskapen 1
2616 Gemenskapens 3
2617 Gemenskapsinitiativet 5
2618 Gemenskapsrätten 1
2619 Gemenskapsåtgärder 2
2620 Genast 1
2621 Gender 1
2622 Generaldirektorat 1
2623 Generaldirektoraten 1
2624 Generaldirektoratet 9
2625 Generaldirektören 1
2626 Generellt 1
2627 Genetiskt 2
2628 Genialiskt 1
2629 Genom 70
2630 Genomförande 1
2631 Genomförandet 4
2632 Genomsnittet 1
2633 Gentila 1
2634 Genua 1
2635 Genève 16
2636 Genèvekonventionen 7
2637 Genèvekonventionens 2
2638 Genèvekonventionerna 1
2639 Genèvemötet 1
2640 George 18
2641 Georges 1
2642 Georgievski 1
2643 Ger 2
2644 Geremek 2
2645 Geresta 1
2646 Getsemane 1
2647 Ghana 1
2648 Ghilardotti 1
2649 Ghoulen 1
2650 Gibraltar 1
2651 Gil-Delgado 1
2652 Gil-Robles 2
2653 Gilderoy 1
2654 Gillig 1
2655 Ginens 1
2656 Ginny 3
2657 Gino 1
2658 Giorgos 5
2659 Gissa 1
2660 Givet 1
2661 Givetvis 6
2662 Gjort 1
2663 Glansen 1
2664 Glase 1
2665 Glasgow 2
2666 Gligorov 1
2667 Global 1
2668 Globaliseringen 5
2669 Globaliseringens 1
2670 Glöm 1
2671 God 1
2672 Goddag 1
2673 Godkännandet 1
2674 Godspeed 1
2675 Goebbels 5
2676 Golan 6
2677 Golanhöjden 1
2678 Golanhöjderna 3
2679 Golden 1
2680 Golfströmmen 3
2681 Golgatavandring 1
2682 Gollnisch 2
2683 Gomes 1
2684 Gong-rörelsen 1
2685 González 2
2686 Goodwill 1
2687 Goodyear 14
2688 Gordon 1
2689 Gorka 1
2690 Gorostiaga 2
2691 Gorsel 3
2692 Gott 2
2693 Gouges 1
2694 Graal 1
2695 Graca 3
2696 Graco-affärerna 1
2697 Graefe 9
2698 Graham 1
2699 Gran 1
2700 Granada 1
2701 Grand 1
2702 Granger 5
2703 Grangers 1
2704 Granskningarna 1
2705 Granskningen 1
2706 Grants 1
2707 Grappakrigen 1
2708 Grattis 2
2709 Gratulerar 1
2710 Gravesend 1
2711 Gray's 1
2712 Graça 5
2713 Great 1
2714 Green 2
2715 Greenspan 1
2716 Greenwich 1
2717 Grekland 42
2718 Greklands 5
2719 Gringotts 4
2720 Grossetête 4
2721 Grosstête 1
2722 Grottor 1
2723 Group 1
2724 Grova 1
2725 Grozny 3
2726 Grunden 4
2727 Grunderna 1
2728 Grundläggande 1
2729 Gruppen 43
2730 Gruppering 1
2731 Grupperna 1
2732 Gruppnivåegenskaper 1
2733 Gruson 1
2734 Gryffindor 1
2735 Grädde 1
2736 Gränsarbetare 1
2737 Gränser 2
2738 Grått 1
2739 Gröna 3
2740 Gröner 2
2741 Grönitz 1
2742 Guatemala 1
2743 Gud 11
2744 Guds 3
2745 Guigou 1
2746 Guld- 1
2747 Guldsökare 1
2748 Gulfkriget 1
2749 Gulfområdet 1
2750 Gusp 1
2751 Guterres 11
2752 Guterrez 1
2753 Gutierres 1
2754 Gutíerrez 2
2755 Gwenzi 1
2756 Gwenzis 1
2757 Gyllenroy 3
2758 Gällande 1
2759 Gärna 1
2760 Gå 2
2761 Gång 2
2762 Går 1
2763 Gör 3
2764 Göra 1
2765 Göteborg 1
2766 Günther 1
2767 H-0002/99 1
2768 H-0006/00 1
2769 H-0020/00 1
2770 H-0021/00 1
2771 H-0022/00 1
2772 H-0024/00 1
2773 H-0025/00 1
2774 H-0026/00 1
2775 H-0027/00 1
2776 H-0028/00 1
2777 H-0029/00 1
2778 H-0031/00 1
2779 H-0035/00 1
2780 H-0036/00 1
2781 H-0040/00 1
2782 H-0041/00 1
2783 H-0042/00 1
2784 H-0044/00 1
2785 H-0045/00 1
2786 H-0045/99 1
2787 H-0049/00 1
2788 H-0052/00 1
2789 H-0053/00 1
2790 H-0057/00 1
2791 H-0095/00 1
2792 H-0117/00 1
2793 H-0122/00 1
2794 H-0209/99 1
2795 H-0218/97 1
2796 H-0237/97 1
2797 H-0778/99 1
2798 H-0780/99 1
2799 H-0781/99 1
2800 H-0782/99 1
2801 H-0785/99 1
2802 H-0786/99 1
2803 H-0788/99 1
2804 H-0791/99 1
2805 H-0793/99 1
2806 H-0795/99 1
2807 H-0796/99 1
2808 H-0798/99 1
2809 H-0801/99 1
2810 H-0805/99 1
2811 H-0807/99 1
2812 H-0808/99 1
2813 H-0813/99 1
2814 H-0817/99 1
2815 H-0819/99 1
2816 H-0829/99 1
2817 H. 1
2818 H.C. 1
2819 HELP 1
2820 HON 1
2821 HOTREC 1
2822 HTML 7
2823 HTML-formatet 1
2824 HTML-kod 1
2825 Ha 1
2826 Haag 3
2827 Haarder 5
2828 Habana 1
2829 Habitat 1
2830 Hade 4
2831 Hadera 1
2832 Hagrid 7
2833 Hague 1
2834 Haider 26
2835 Haiderpolitiken 1
2836 Haiders 24
2837 Haifa 1
2838 Hain 1
2839 Hainaut 1
2840 Halonen 1
2841 Halva 1
2842 Hamburg 2
2843 Hamilton 1
2844 Hamna 1
2845 Hamnarna 1
2846 Hamnens 1
2847 Han 378
2848 Handeln 1
2849 Handelsavtal 1
2850 Handelsavtalet 1
2851 Handicap 1
2852 Handikappades 1
2853 Handikapporganisationer 1
2854 Handlingen 1
2855 Handlingskraften 1
2856 Hangarfartyget 1
2857 Hannas 1
2858 Hans 28
2859 Hanteringen 1
2860 Har 33
2861 Harbour 2
2862 Harbours 1
2863 Harmoniseringsbyrån 1
2864 Harold 1
2865 Harpoon 1
2866 Harry 147
2867 Harrys 18
2868 Harvey 1
2869 Harveys 1
2870 Harwich 1
2871 Hatzidakis 3
2872 Hatzidakisbetänkandet 1
2873 Haug 1
2874 Hautala 4
2875 Havel 10
2876 Havels 2
2877 Haven 1
2878 Havet 1
2879 Havsprodukternas 1
2880 Havsvärlden 1
2881 Heathrow 2
2882 Heaton-Harris 1
2883 Hebreiska 1
2884 Hebriderna 1
2885 Hebron- 1
2886 Hecke 3
2887 Heckes 2
2888 Hedge 1
2889 Hedkvist 1
2890 Hedwig 5
2891 Hedwig's 1
2892 Hedwigs 2
2893 Hefaistos 1
2894 Heidi 1
2895 Heights 1
2896 Heinz 1
2897 Hej 2
2898 Hela 15
2899 Helighet 1
2900 Helmkom-avtalet 1
2901 Helms-Burton 1
2902 Help 1
2903 Helsingfors 52
2904 Helsingfors-besluten 1
2905 Helsingforskonventionen 1
2906 Helsingforsmandatet 1
2907 Helsingforsmötet 2
2908 Helsingforstoppmötet 1
2909 Helt 8
2910 Hemliga 1
2911 Hemma 1
2912 Hennes 13
2913 Henry 3
2914 Hereford 1
2915 Herman 2
2916 Hermes 1
2917 Hermione 10
2918 Hernandez 1
2919 Hernando 1
2920 Hernández 1
2921 Herr 967
2922 Herre 1
2923 Herregud 1
2924 Herritarrok 2
2925 Hertfordshire 1
2926 Hicks 1
2927 Hilton 1
2928 Himalaya 1
2929 Himalayabergen 1
2930 Hind 1
2931 Hindenburg 1
2932 Hinken 1
2933 Hinner 1
2934 Historia 1
2935 Historien 6
2936 Hit 4
2937 Hitler 11
2938 Hitler-regimen 1
2939 Hitlers 1
2940 Hittar 1
2941 Hittills 8
2942 Hjalmar 9
2943 Hjälp 3
2944 Hoechst 1
2945 Hogwarts 16
2946 Holland 3
2947 Hollywoodfilmer 1
2948 Holzmann 1
2949 Holzmann-gruppen 1
2950 Hon 91
2951 Honduras 2
2952 Hong 1
2953 Hongkong 4
2954 Hoogoven 1
2955 Hopkerk 1
2956 Hoppet 2
2957 Horizon 2
2958 Horst 1
2959 Hos 1
2960 Hotel 5
2961 Hotelsemönstret 1
2962 Hoti 1
2963 House 2
2964 Hover 1
2965 Howard 1
2966 Howittsbetänkandet 1
2967 Hubert 1
2968 Hudghton 8
2969 Hudghtons 1
2970 Hudsonfloden 1
2971 Hugg 1
2972 Hughes 1
2973 Huhne 5
2974 Huj 4
2975 Hulten 12
2976 Hultenbetänkandet 4
2977 Hultens 3
2978 Hulthen 4
2979 Hulthens 2
2980 Human 1
2981 Hun 1
2982 Hundratals 1
2983 Hungersnöd 1
2984 Hur 119
2985 Hurdana 1
2986 Huruvida 3
2987 Huset 1
2988 Hustrun 2
2989 Huvudaktörerna 1
2990 Huvudansvaret 1
2991 Huvudbudskapet 1
2992 Huvuddelen 1
2993 Huvudfrågorna 1
2994 Huvudlinjen 1
2995 Huvudmålet 1
2996 Huvudmålsättningen 1
2997 Huvudproblemet 1
2998 Huvudregeln 1
2999 Huvudsaken 3
3000 Hyckleri 1
3001 Hypertext 1
3002 Häkkinens 1
3003 Häktningsorder 1
3004 Hälften 1
3005 Händelsen 1
3006 Händelser 1
3007 Händelserna 3
3008 Hängde 1
3009 Hänsch 2
3010 Hänsyn 3
3011 Här 86
3012 Härav 2
3013 Härigenom 1
3014 Härmed 6
3015 Härom 1
3016 Häromdagen 1
3017 Hästen 2
3018 Håll 3
3019 Hållbar 2
3020 Håller 1
3021 Hår 1
3022 Hög 3
3023 Höga 1
3024 Högaktningsfullt 1
3025 Höge 1
3026 Högerextremism 1
3027 Högnivågruppen 2
3028 Högre 1
3029 Högst 1
3030 Högvärdighet 1
3031 Höjden 1
3032 Hör 1
3033 I 907
3034 I-programmet 2
3035 I. 1
3036 IBM 1
3037 ICCAT 6
3038 ICCAT:s 2
3039 ICES 1
3040 ICES-zon 1
3041 ICES-zonen 1
3042 ICES-zonerna 1
3043 ICT-företag 1
3044 ID 1
3045 IDEA-åldern 1
3046 IFOP 1
3047 IGC 4
3048 II 28
3049 II-programmet 4
3050 III 26
3051 III- 1
3052 III-gränser 1
3053 III-initiativet 1
3054 III-programmet 2
3055 IIIA 1
3056 IIIC 2
3057 ILA 21
3058 ILO 2
3059 IMF 1
3060 IMO 2
3061 IMO:s 1
3062 INTE 1
3063 INTERREG 2
3064 INTERREG-initiativ 1
3065 IOPCF 2
3066 IOPCF:s 1
3067 IRA 1
3068 ISA 1
3069 ISD 1
3070 ISPA-instrumentet 1
3071 IT 9
3072 IT-branschen 1
3073 IT-fattiga 1
3074 IT-infrastruktur 2
3075 IT-rika 1
3076 IT-utvecklingen 1
3077 ITALIENSKA 1
3078 IV 5
3079 IX 2
3080 Ibland 9
3081 Icke 6
3082 Icke-statliga 1
3083 Identifiera 1
3084 Idén 3
3085 Igal 1
3086 Igår 1
3087 Ihållande 1
3088 Ikväll 1
3089 Ile-de-France 1
3090 Ilisu- 1
3091 Ilisudammen 4
3092 Illa 1
3093 Illegalt 1
3094 Ilsket 1
3095 Imbeni 3
3096 Immigrationen 1
3097 Immobile 1
3098 Importera 4
3099 Inbillar 1
3100 Inbjudningarna 1
3101 Inbördes 1
3102 Independence 1
3103 Indien 6
3104 Indiens 1
3105 Indikatorerna 1
3106 Indirekt 1
3107 Indiska 1
3108 Indonesien 11
3109 Industriella 1
3110 Industrin 1
3111 Industrins 1
3112 Infektiös 1
3113 Information 2
3114 Informationen 2
3115 Informationscentren 1
3116 Informationssamhället 1
3117 Infödingsmattor 1
3118 Inför 10
3119 Införandet 4
3120 Inga 8
3121 Ingen 30
3122 Ingenstans 2
3123 Ingenting 5
3124 Inger 1
3125 Inget 9
3126 Ingetdera 1
3127 Inglewood 1
3128 Inglewoods 1
3129 Ingusjien 1
3130 Initiativ 1
3131 Initiativet 6
3132 Initiativets 1
3133 Inklusive 1
3134 Inkomstklyftan 1
3135 Inlåst 1
3136 Inlåsta 1
3137 Inn 1
3138 Innan 22
3139 Innebär 1
3140 Innebörden 1
3141 Innehållet 1
3142 Innehållsmässigt 1
3143 Innovation 1
3144 Inom 30
3145 Inre 2
3146 Inresan 1
3147 Inriktning 1
3148 Inrättandet 1
3149 Insamling 1
3150 Insatserna 2
3151 Insatsstyrkan 1
3152 Inskränkningarna 1
3153 Insolvens 1
3154 Insolvensförfaranden 1
3155 Installera 1
3156 Institute 1
3157 Institutionellt 1
3158 Instrumenten 2
3159 Inte 70
3160 Integra 2
3161 Integritet 1
3162 Intellectual 2
3163 Intern 1
3164 International 7
3165 Internationell 2
3166 Internationella 25
3167 Internet 42
3168 Internet-ekonomins 1
3169 Internetrevolutionen 2
3170 Internetrevolutionens 1
3171 Interreg 71
3172 Interreg- 1
3173 Interreg-anslag 1
3174 Interreg-anslagen 1
3175 Interreg-initiativ 1
3176 Interreg-initiativet 9
3177 Interreg-programmen 1
3178 Interreg-programmet 2
3179 Interreg-riktlinjer 1
3180 Interreg-ärendena 1
3181 Interregs 4
3182 Interventionspriser 1
3183 Intill 2
3184 Intressant 2
3185 Invandrarna 1
3186 Investeringar 2
3187 Investeringsnivåerna 1
3188 Investments 1
3189 Ionescu 1
3190 Irak 5
3191 Iraks 1
3192 Iran 3
3193 Irans 1
3194 Irland 52
3195 Irlands 2
3196 Irländska 7
3197 Isabel 3
3198 Island 1
3199 Isler 2
3200 Ismail 1
3201 Isoza-floden 1
3202 Ispa 1
3203 Ispa- 1
3204 Ispar 1
3205 Israel 84
3206 Israel-Syrienfrågan 1
3207 Israeliska 1
3208 Israelkritik 1
3209 Israels 18
3210 Istanbul 1
3211 Istället 5
3212 Italien 41
3213 Italiens 1
3214 Ivanov 1
3215 Izquierdo 1
3216 J 3
3217 JAG 1
3218 Ja 64
3219 Ja-så-är-vi-här-igen-leende 1
3220 Jackson 2
3221 Jacob 2
3222 Jacques 8
3223 Jaffa 2
3224 Jag 2966
3225 Jaga 1
3226 Jaha 2
3227 Jakov 1
3228 Jalta 1
3229 Jamaica 2
3230 Jamen 3
3231 James 6
3232 Jan 3
3233 Jan-Kees 1
3234 Jan-feb 1
3235 Japan 9
3236 Jarzembowski 3
3237 Jason 2
3238 Jaså 5
3239 Javette-Le 1
3240 Javier 9
3241 Jean 5
3242 Jean-Claude 2
3243 Jean-Olivier 1
3244 Jefferson 1
3245 Jens-Peter 1
3246 Jeremia 1
3247 Jersey 2
3248 Jerusalem 13
3249 Jerusalems 4
3250 Jesus 2
3251 Jet 1
3252 Jo 8
3253 Jo-Ann 2
3254 Joakim 1
3255 Joaquim 1
3256 Joaquín 1
3257 Jobert 1
3258 Jobs 2
3259 Jodå 1
3260 Johan 1
3261 Johannes' 1
3262 John 17
3263 Jojon 2
3264 Jomän 1
3265 Jonas 2
3266 Jonckheer 9
3267 Jonckheerbetänkandet 3
3268 Jonckheers 3
3269 Jord 1
3270 Jordan 1
3271 Jordanien 1
3272 Jordanierna 1
3273 Jordans 1
3274 Jordbruk 2
3275 Jordbrukande 1
3276 Jordbruket 3
3277 Jordbruksekonomin 1
3278 Jordbruksministeriet 1
3279 Jorge 3
3280 Josafats 1
3281 Joseph 1
3282 Jospin 3
3283 José 2
3284 Journal 1
3285 Journalisten 1
3286 Journalister 2
3287 Journalists 1
3288 Jove 5
3289 Jovisst 1
3290 Joyces 1
3291 Ju 6
3292 Judarna 1
3293 Judeens 1
3294 Judegrabbens 1
3295 Judismen 1
3296 Jugoslavien 32
3297 Jugoslaviens 7
3298 Juncker 1
3299 Jung 1
3300 Junker 1
3301 Junkers 1
3302 Juridisk 1
3303 Just 36
3304 Justering 7
3305 Justeringen 1
3306 Jämförelse 1
3307 Jämfört 4
3308 Jämställdhet 2
3309 Jämställdheten 1
3310 Jämställdhetsaspekter 1
3311 Jörg 18
3312 Jösses 2
3313 Júcar 2
3314 KFOR 1
3315 KLM 1
3316 KOM(1997 1
3317 KOM(1998 5
3318 KOM(1999 21
3319 KOM(1999)0003 2
3320 KOM(1999)0598 1
3321 KOM(98)0662 1
3322 KOM(99)0598 1
3323 Kabila 1
3324 Kabul 1
3325 Kackerlackor 1
3326 Kafferast 1
3327 Kafor 1
3328 Kairo 2
3329 Kaleidoskop 2
3330 Kalejdoskop 1
3331 Kambodja 14
3332 Kambodjas 1
3333 Kammaren 5
3334 Kampen 1
3335 Kan 53
3336 Kanada 6
3337 Kanarieöarna 2
3338 Kandalprovinsen 1
3339 Kandidatländerna 1
3340 Kandidatländernas 1
3341 Kano 1
3342 Kanske 23
3343 Kantabrien 3
3344 Kapital- 1
3345 Kaptenen 1
3346 Karamanous 1
3347 Karas 4
3348 Karelen 1
3349 Karibien 5
3350 Karin 1
3351 Karl 6
3352 Karl-Heinz 2
3353 Karlsruhe 2
3354 Kartellamt 1
3355 Kartellförbudet 1
3356 Kaspiska 1
3357 Katalonien 1
3358 Katastrofen 1
3359 Katastrofer 1
3360 Kategorifältområde 1
3361 Katharine 1
3362 Katiforis 26
3363 Katiforisbetänkandet 2
3364 Kattflatan 1
3365 Kaufmann 1
3366 Kaukasus 4
3367 Kauppi 2
3368 Kazakstan 1
3369 Kedourie 3
3370 Kedouries 1
3371 Kejsarens 1
3372 Kellett-Bowman 1
3373 Kemikalier 1
3374 Kennedy 1
3375 Kensington 1
3376 Kente 2
3377 Kenyatta 1
3378 Kermit 1
3379 Kfor 1
3380 Kfor-styrkan 1
3381 Kfor-styrkorna 1
3382 Kfor-trupperna 1
3383 Khartum 1
3384 Khatami 2
3385 Kina 45
3386 Kinapolitik 1
3387 Kinas 4
3388 Kindermann 3
3389 King 1
3390 Kinnock 29
3391 Kinnocks 5
3392 Kippur 1
3393 Kirgizistan 5
3394 Kissinger 2
3395 Kit 1
3396 Kjolarna 1
3397 Klart 1
3398 Klicka 1
3399 Klimas 1
3400 Klippan 1
3401 Klistra 1
3402 Klockan 6
3403 Knappt 1
3404 Knörr 7
3405 Koch 15
3406 Kochs 1
3407 Kocken 1
3408 Kod 1
3409 Kodaks 1
3410 Koden 1
3411 Kofi 1
3412 Kohl 1
3413 Kohoutek 1
3414 Kollega 1
3415 Kollegan 3
3416 Kolleger 3
3417 Kollektiva 1
3418 Kom 7
3419 Kombinera 1
3420 Kommandot 1
3421 Kommer 34
3422 Kommissarie 1
3423 Kommissionen 202
3424 Kommissionens 62
3425 Kommissionsledamöterna 1
3426 Kommissionär 22
3427 Kommissionären 9
3428 Kommissionärerna 1
3429 Kommittologi 1
3430 Kommittéförfarande 2
3431 Kommitténs 1
3432 Kommuner 1
3433 Kommunerna 1
3434 Kompletterande 1
3435 Kompromissformuleringar 1
3436 Koncentrationen 1
3437 Konceptet 2
3438 Konflikten 2
3439 Kong 1
3440 Kongo 7
3441 Kongressen 1
3442 Kongs 1
3443 Konkret 1
3444 Konkreta 1
3445 Konkurrens 3
3446 Konkurrensen 6
3447 Konkurrenspolitik 1
3448 Konkurrenspolitiken 4
3449 Konkurrensprincipen 2
3450 Konrad 1
3451 Konsekvenserna 3
3452 Konstigt 1
3453 Konsumenten 1
3454 Konsumenterna 4
3455 Konsumentpolitiken 1
3456 Kontoren 1
3457 Kontroll 1
3458 Kontroller 4
3459 Kontrollfunktionen 1
3460 Kontrollförfarandet 1
3461 Kontrollnamn 1
3462 Kontrollpanel 1
3463 Kontrollstöd 1
3464 Konventionen 4
3465 Konventioner 1
3466 Konvertera 1
3467 Kopiera 3
3468 Kopplat 1
3469 Korea 3
3470 Korrekt 1
3471 Korridorerna 1
3472 Kors 1
3473 Korsfrågor 1
3474 Kort 11
3475 Kortfattat 2
3476 Koschermat 1
3477 Kososvokonflikten 1
3478 Kosova 1
3479 Kosovo 176
3480 Kosovoalbanerna 1
3481 Kosovofrågan 1
3482 Kosovoinsatser 1
3483 Kosovokonflikten 3
3484 Kosovokriget 2
3485 Kosovokrigets 1
3486 Kosovoproblemet 1
3487 Kosovos 17
3488 Kostnaden 1
3489 Kostnaderna 5
3490 Kotka 1
3491 Kouchener 1
3492 Kouchner 14
3493 Kouchners 9
3494 Koushner 1
3495 Koushners 2
3496 Kraftiga 1
3497 Krajina 1
3498 Krav 1
3499 Kraven 1
3500 Kravet 2
3501 Kreml 2
3502 Kriget 3
3503 Krigsherrar 1
3504 Kriterier 1
3505 Kroatien 6
3506 Kronos 1
3507 Kroppen 1
3508 Kuba 22
3509 Kubas 6
3510 Kuckelkorn 1
3511 Kultur 20
3512 Kulturell 3
3513 Kulturellt 1
3514 Kulturen 1
3515 Kumar 1
3516 Kunde 1
3517 Kunder 2
3518 Kundorder 1
3519 Kungliga 1
3520 Kunskapssamhället 1
3521 Kurti 1
3522 Kurtz 10
3523 Kusligt 1
3524 Kuwait 1
3525 Kv3 1
3526 Kvalitet 2
3527 Kvalitén 1
3528 Kvantifierade 1
3529 Kvartal 1
3530 Kvestorerna 1
3531 Kvicksilver 1
3532 Kvinnan 2
3533 Kvinnor 22
3534 Kvinnorna 7
3535 Kvinnornas 4
3536 Kvinnors 2
3537 Kvotering 1
3538 Kväkareuropa 1
3539 Kyi 1
3540 Kyoto 6
3541 Kyoto-protokollet 1
3542 Kyotoprocesserna 1
3543 Kyotoprotokollet 2
3544 Kyotos 1
3545 Kypare 1
3546 Kyrkans 1
3547 Känner 4
3548 Känsliga 1
3549 Kära 18
3550 Käraste 1
3551 Käre 1
3552 Kärnan 1
3553 Kärnkraftverk 1
3554 Kärnkraftverket 1
3555 Kärnten 3
3556 Köhler 1
3557 Köket 1
3558 Köln 7
3559 Kölnprocessen 2
3560 Kön 1
3561 Köp 1
3562 Köpenhamn 4
3563 L 1
3564 LEVE 1
3565 LIMIT 1
3566 LOCKMAN 1
3567 LTCM 1
3568 La 8
3569 Laan 2
3570 Laans 5
3571 Labourregeringens 1
3572 Labours 1
3573 Labrador 1
3574 Lagkatalogen 1
3575 Lagstiftningen 1
3576 Lama 5
3577 Lamas 2
3578 Lambala 1
3579 Lambalas 1
3580 Lancker 3
3581 Land 1
3582 Landaburu 1
3583 Landet 4
3584 Landis 1
3585 Landsbygden 1
3586 Landsbygdens 1
3587 Landsbygdsområdena 1
3588 Lange 12
3589 Langen 13
3590 Langenbetänkandet 1
3591 Langens 3
3592 Langer 2
3593 Langes 1
3594 Language 6
3595 Lanka 3
3596 Lannoye 4
3597 Lannoyes 1
3598 Lappland 3
3599 Lapus 1
3600 Larcher 1
3601 Lastbilen 1
3602 Lastbilstrafiken 1
3603 Lasten 1
3604 Latina 2
3605 Latinamerika 1
3606 Laurent 1
3607 Le 6
3608 Leader 47
3609 Leader+ 25
3610 Leader+-initiativen 1
3611 Leader+-programmen 1
3612 Leader+-programmet 6
3613 Leader-initiativet 3
3614 Leader-programmen 1
3615 Leader-programmens 1
3616 Leader-programmet 4
3617 Leader-projekten 1
3618 Leader-stödområdena 1
3619 Lechner 2
3620 Leclerc 1
3621 Ledamot 4
3622 Ledamoten 7
3623 Ledamotens 1
3624 Ledamöter 4
3625 Ledamöterna 2
3626 Ledare 1
3627 Ledley 1
3628 Ledningen 1
3629 Lee 1
3630 Leendet 1
3631 Legenden 2
3632 Leinemanns 2
3633 Leinen 7
3634 Leinens 1
3635 Leinster 1
3636 Leinsters 1
3637 Leon 1
3638 Leonardo 1
3639 Leone 1
3640 Leoni 1
3641 Lepers 1
3642 Lepos 1
3643 Lesotho 1
3644 Lettland 1
3645 Lev 1
3646 Levande 1
3647 Levante 1
3648 Levantines 2
3649 Libanon 6
3650 Liberal 2
3651 Liberaliseringen 1
3652 Liberty 2
3653 Libyens 1
3654 License 1
3655 Lider 1
3656 Lieneman 1
3657 Lienemann 19
3658 Lienemannbetänkandet 1
3659 Lienemanns 9
3660 Lienemannsbetänkandet 1
3661 Life 52
3662 Life-Miljö 1
3663 Life-Natur 1
3664 Life-Tredje 1
3665 Life-förordningen 1
3666 Life-instrumentet 1
3667 Life-miljö 1
3668 Life-natur 1
3669 Life-programmen 1
3670 Life-programmet 2
3671 Life-programmets 1
3672 Life-projekt 1
3673 Life-projektets 1
3674 Life:s 2
3675 Lifes 1
3676 Liikanen 14
3677 Lika 1
3678 Likadant 1
3679 Likafullt 2
3680 Likaså 6
3681 Like 1
3682 Liknande 1
3683 Likriktning 1
3684 Liksom 18
3685 Likväl 4
3686 Lille 1
3687 Lillehammer-rapporten 1
3688 Limpopodalen 1
3689 Lindgren 2
3690 Linds 1
3691 Link 1
3692 Links 1
3693 Lipietz 1
3694 Lissabon 83
3695 Lissabon-initiativ 1
3696 Lissabonmötet 4
3697 Listorna 1
3698 Litauen 3
3699 Lite 1
3700 Litteraturen 1
3701 Little 1
3702 Liverpool 3
3703 Livet 1
3704 Livliga 9
3705 Livsmedelssäkerhet 2
3706 Livsmedelssäkerheten 2
3707 Livsmedelssäkerhetsmyndigheten 1
3708 Livsmedelssäkerhetsprogram 1
3709 Livsmedelsäkerhet 1
3710 Ljuden 1
3711 Ljug 1
3712 Ljuspunkterna 1
3713 Lloyds 1
3714 Lockhart 1
3715 Lockman 3
3716 Lockmans 1
3717 Logiskt 1
3718 Loi 1
3719 Loire 1
3720 Loire-Atlantique 2
3721 Lokala 1
3722 Lomas 1
3723 Lomé 3
3724 Loméavtal 1
3725 Loméavtalens 1
3726 Loméavtalet 2
3727 Lomékonvention 1
3728 Lomékonventionen 18
3729 Lomékonventionens 3
3730 Lomékonventionerna 1
3731 Loméländerna 1
3732 Lomémodellen 1
3733 Loméramen 1
3734 Lomésamarbetet 1
3735 Loméuppgörelse 1
3736 London 17
3737 Lord 4
3738 Lorenzettis 1
3739 Lorosae 1
3740 Lorraine 2
3741 Lothar 3
3742 Louis 4
3743 Lousewies 1
3744 Louth 1
3745 Loyola 2
3746 Lucas 6
3747 Lucius 1
3748 Luften 3
3749 Lugard 1
3750 Luis 2
3751 Lukten 1
3752 Lulling 2
3753 Luncheonette 1
3754 Lund 2
3755 Luren 1
3756 Lutte 1
3757 Luxemburg 21
3758 Luxemburgprocess 3
3759 Luxemburgprocessen 6
3760 Luxemburgprocessens 1
3761 Luxemburgs 1
3762 Luxemburgstrategin 1
3763 Lycka 1
3764 Lyckas 1
3765 Lyckligt- 1
3766 Lyckligtvis 4
3767 Lydda 1
3768 Lyncharna 1
3769 Lynne 2
3770 Lynnes 2
3771 Lyon 1
3772 Lyssna 1
3773 LÄRT 1
3774 Läge 1
3775 Läget 3
3776 Lägg 7
3777 Lägga 2
3778 Lägre 1
3779 Lämna 1
3780 Lämnade 1
3781 Lämplig 1
3782 Lämpliga 1
3783 Lämpligt 1
3784 Länder 2
3785 Längs 1
3786 Länka 2
3787 Lärande 1
3788 Läs 3
3789 Lån 1
3790 Långrandigt 1
3791 Långsamheten 1
3792 Långt 1
3793 Låt 150
3794 Lönsamhet 1
3795 Lösningarna 1
3796 Lösningen 3
3797 Lööw 2
3798 Lübeck 1
3799 MAGISK 1
3800 MARPOL 1
3801 MATEN 1
3802 MPLA 2
3803 MSDN 1
3804 MSF 1
3805 MUTE 1
3806 Maaaaaammma 1
3807 Maastricht 4
3808 Maastrichtfördraget 8
3809 Maastrichtkonferensen 1
3810 Maastrichtkriterierna 2
3811 Maaten 3
3812 MacCormick 6
3813 Macao 2
3814 Mace 1
3815 Machie 1
3816 Mad 1
3817 Madagaskar 2
3818 Madeira 3
3819 Madison 2
3820 Madrid 4
3821 Madrid- 1
3822 Maes 6
3823 Mafalda 1
3824 Maghreb 1
3825 Maghrebländerna 1
3826 Maij-Weggen 4
3827 Maij-Weggens 1
3828 Mainstreaming 1
3829 Majestäts 2
3830 Major 1
3831 Majoriteten 3
3832 Makedonien 66
3833 Makedoniens 5
3834 Makten 1
3835 Maktproblem 1
3836 Malenga 1
3837 Malfoy 14
3838 Malfoys 1
3839 Mallorca 1
3840 Malmström 3
3841 Malone 1
3842 Malta 42
3843 Maltas 4
3844 Mamma 2
3845 Mamère 1
3846 Man 196
3847 Managing 1
3848 Manchester 2
3849 Mandela 1
3850 Mandelstam 2
3851 Manes 1
3852 Manhattan 1
3853 Mannen 7
3854 Mansons 1
3855 Manuel 1
3856 Manyema 1
3857 Mappen 1
3858 Maputo 1
3859 Mar-Apr 1
3860 Marches 1
3861 Mare 1
3862 Margarin 1
3863 Marginaliseringen 1
3864 Margot 12
3865 Maria 2
3866 Marie 1
3867 Marie-Noëlle 2
3868 Marindepartementet 1
3869 Marinho 5
3870 Marinhos 1
3871 Mario 2
3872 Maritain 1
3873 Markera 1
3874 Marknaden 5
3875 Marknadsverkan 1
3876 Markov 4
3877 Markup 2
3878 Marlow 4
3879 Marlows 1
3880 Marocko 7
3881 Marpol-fördraget 1
3882 Marpolkonventionen 2
3883 Marques 1
3884 Marseille 1
3885 Marset 1
3886 Marshallplan 1
3887 Marshallplanen 1
3888 Marshallplaner 1
3889 Martin 5
3890 Martinez 2
3891 Martini 1
3892 Martín 4
3893 Martíns 1
3894 Masker 1
3895 Mason 5
3896 Masons 1
3897 Massor 1
3898 Matematiker 1
3899 Maten 1
3900 Mathieu 1
3901 Matisse 1
3902 Matrovica 1
3903 Matrovicas 1
3904 Maurice 1
3905 Max 2
3906 Maximalt 1
3907 Maximiåldern 1
3908 McCarthy 7
3909 McCartin 1
3910 McGowan 1
3911 McKenna 2
3912 McNally 3
3913 McNallybetänkandet 1
3914 McNallys 1
3915 Meat 1
3916 Mebeki 1
3917 Med 153
3918 Meda 7
3919 Meda-programmet 2
3920 Medan 28
3921 Medbeslutande 1
3922 Medborgare 2
3923 Medborgaren 1
3924 Medborgarna 7
3925 Medborgarnas 1
3926 Meddelande 1
3927 Medel 1
3928 Medelhavet 22
3929 Medelhavets 5
3930 Medelhavshamnar 2
3931 Medelhavsländer 1
3932 Medelhavsländerna 5
3933 Medelhavsområdet 8
3934 Medelhavsområdets 1
3935 Medelhavsregionen 2
3936 Medelhavstonfisken 1
3937 Medellängd 1
3938 Medger 1
3939 Medicinen 1
3940 Medina 5
3941 Medlemsstaterna 13
3942 Medlemsstaternas 3
3943 Medresenärerna 1
3944 Medvetandet 1
3945 Meijer 1
3946 Mekanisk 1
3947 Mellan 5
3948 Mellanöstern 45
3949 Mellanösternfreden 1
3950 Mellanösternkampen 1
3951 Mellanösternpolitik 1
3952 Mellanösterns 2
3953 Melville 2
3954 Melvilles 1
3955 Memoirs 1
3956 Men 627
3957 Menar 3
3958 Meningen 2
3959 Mentaliteten 1
3960 Menéndez 1
3961 Mer 19
3962 Merseybeat 1
3963 Messias 1
3964 Messieurs 1
3965 Mest 1
3966 Metallräcket 1
3967 Metis 3
3968 Mets 5
3969 Mexico 1
3970 Mexiko 3
3971 Michel 5
3972 Michelin 4
3973 Michelin-koncernen 1
3974 Michiel 1
3975 Microsoft 37
3976 Middelhoek 1
3977 Midlands 2
3978 Miert 1
3979 Miggs 1
3980 Mika 1
3981 Milano 1
3982 Milano-området 1
3983 Miles 1
3984 Militär 1
3985 Miljoner 1
3986 Miljöaspekterna 1
3987 Miljöinstitutioner 1
3988 Miljökatastrof 1
3989 Miljökatastrofen 1
3990 Miljökatastroferna 1
3991 Miljömässigt 1
3992 Miljön 2
3993 Miljöproblem 1
3994 Miljöproblemen 1
3995 Miljösituationen 1
3996 Miljövariabeln 1
3997 Millennierundan 1
3998 Millennium 3
3999 Miller 3
4000 Milosevic 11
4001 Milosevic-regimen 1
4002 Milosevicregimen 1
4003 Milosevics 6
4004 Min 118
4005 Mina 37
4006 Minchah-bön 1
4007 Mindre 2
4008 Minimiregler 1
4009 Minimistorleken 1
4010 Minister 2
4011 Ministeriet 3
4012 Ministern 2
4013 Ministerrådet 1
4014 Minnen 1
4015 Minnesota 1
4016 Minns 2
4017 Minoriteter 1
4018 Minsk 1
4019 Minskar 1
4020 Minskningen 1
4021 Minst 1
4022 Minsta 1
4023 Minuc 1
4024 Mira 2
4025 Mirakel 1
4026 Miranda 1
4027 Mishkenot 1
4028 Mississippi 2
4029 Mister 2
4030 Mitrovic 1
4031 Mitrovica 17
4032 Mitt 20
4033 Mittemot 1
4034 Mitterrand 1
4035 Mitterrands 1
4036 Moabs 1
4037 Mobiliseringen 1
4038 Moby 1
4039 Moder 2
4040 Modern 1
4041 Modernare 1
4042 Modernisering 1
4043 Modrow 1
4044 Mohieddin 1
4045 Moldavien 1
4046 Mollar 2
4047 Molly 3
4048 Moloksdyrkarna 1
4049 Moluckerna 3
4050 Mom's 1
4051 Monde 5
4052 Mongoliet 2
4053 Monica 1
4054 Monika 2
4055 Monnet 1
4056 Monnets 1
4057 Monsieur 1
4058 Montego 1
4059 Montenegro 2
4060 Monti 28
4061 Monti-paketet 1
4062 Montipaketet 1
4063 Montis 1
4064 Montreal 4
4065 Mor 7
4066 Moral 1
4067 Moratinos 4
4068 Moratorium 1
4069 Morbihan 1
4070 Morbror 5
4071 Morgan 6
4072 Morgantini 5
4073 Morgantinis 1
4074 Morillon 2
4075 Morituri 1
4076 Morse 1
4077 Moseboken 1
4078 Moses 1
4079 Moshe 1
4080 Moskva 3
4081 Moss 1
4082 Moster 4
4083 Mot 27
4084 Motiveringen 1
4085 Motorn 1
4086 Motsättningar 1
4087 Mottagningsanordningar 1
4088 Mount 1
4089 Mountain 4
4090 Moura 8
4091 Mouskouri 1
4092 Mozambique 4
4093 Mozart 1
4094 Moçambique 47
4095 Moçambiques 3
4096 Mr 19
4097 Mrs 20
4098 Msaccess.exe 1
4099 Mugabe 1
4100 Muggle 3
4101 Muggles 4
4102 Mulder 2
4103 Muntorrhet 1
4104 Murcia 1
4105 Murphy 1
4106 Muscardini 1
4107 Muscovy 1
4108 Musik 1
4109 Musiken 1
4110 Musket-skjutning 1
4111 Musselodlingen 1
4112 Mussolinihaka 1
4113 Mweta 30
4114 Mwetas 7
4115 Myanmar 2
4116 Mycket 15
4117 Myller 1
4118 Myndigheten 2
4119 Myndighetens 2
4120 Män 2
4121 Mängden 1
4122 Mängdfunktionerna 1
4123 Människor 6
4124 Människorna 4
4125 Människors 2
4126 Människorättsorganisationen 1
4127 Människorättsorganisationer 1
4128 Människorättspolitiken 1
4129 Mänskliga 9
4130 Mänsklighetens 1
4131 Märkligt 2
4132 Märks 1
4133 Mätare 1
4134 Mätt 1
4135 Må 1
4136 Måhända 1
4137 Målarfärgen 1
4138 Målet 13
4139 Målsättningen 3
4140 Många 36
4141 Månljuset 1
4142 Måste 3
4143 Måtte 2
4144 Méndez 1
4145 Möblerna 1
4146 Möjligen 1
4147 Möjligheten 3
4148 Möjligheter 1
4149 Möjligt 1
4150 Mörkt 1
4151 Möten 1
4152 München 3
4153 Münchens 1
4154 Münchhausen 1
4155 NGL-gruppen 3
4156 NL 7
4157 NT 2
4158 NT-användaren 1
4159 NT-plattform 1
4160 Nagorno-Karabach 2
4161 Namibia 6
4162 Namnet 3
4163 Namnge 1
4164 Nana 1
4165 Nantucket 3
4166 Napoleon 2
4167 Napoleonkrigen 1
4168 Napoleons 1
4169 Napolitano 6
4170 Napolitanos 1
4171 Narcissus 1
4172 Narkotikafrågan 1
4173 Narkotikahandeln 1
4174 Nasdaq 2
4175 Nasdaq- 1
4176 Nassau 3
4177 Nassaumötets 1
4178 Nasser 3
4179 Nassers 3
4180 National 2
4181 Nationaliteter 1
4182 Nationalstaterna 1
4183 Nationella 5
4184 Nationernas 4
4185 Nations 1
4186 Nato 38
4187 Nato-församlingens 1
4188 Nato-länderna 1
4189 Nato-styrkornas 1
4190 Natoaktionen 1
4191 Natobasen 1
4192 Natos 35
4193 Natostyrkor 1
4194 Natostyrkornas 1
4195 Natten 1
4196 Natura 5
4197 Naturliga 1
4198 Naturligtvis 42
4199 Nauvoo 1
4200 Navrozov 2
4201 Neapel 2
4202 Nederländerna 25
4203 Nederländernas 1
4204 Nedläggningen 1
4205 Neil 11
4206 Neils 2
4207 Nej 33
4208 Nellie 1
4209 Ner 1
4210 Nere 1
4211 Nervcentrum 1
4212 Netanyahus 1
4213 Network 1
4214 New 20
4215 Newcastle 1
4216 News 2
4217 Newton 1
4218 Ni 177
4219 Ni-vet-vem 1
4220 Nicaragua 1
4221 Nice 1
4222 Nicholson 1
4223 Nicole 4
4224 Nicosia 1
4225 Nicosias 2
4226 Nielsen 2
4227 Nielsens 1
4228 Nielson 23
4229 Nielsons 3
4230 Nigeria 3
4231 Nikitin 2
4232 Nimbus 1
4233 Nissan 1
4234 Nivån 2
4235 Nja 1
4236 Njaa 1
4237 Nobelpris 1
4238 Nobelpristagare 1
4239 Nog 1
4240 Noggrann 1
4241 Nogueira 4
4242 Noirmoutier 1
4243 Noiz 1
4244 Nord 4
4245 Nord-Pas-de-Calais 1
4246 Nord-Syd 1
4247 Nordafrika 3
4248 Nordatlanten 2
4249 Nordatlantiska 1
4250 Norden 1
4251 Nordeuropa 1
4252 Nordirland 10
4253 Nordirlands 3
4254 Nordisk 7
4255 Norditalien 1
4256 Nordostatlantpakten 1
4257 Nordpolen 1
4258 Nordsjön 3
4259 Nordsjöområdet 1
4260 Norge 13
4261 Norges 1
4262 Normala 1
4263 Normer 1
4264 Norr 1
4265 North 2
4266 Northfield 1
4267 Now 2
4268 Now-projektet 1
4269 Noël 1
4270 Nu 77
4271 Null-värde 1
4272 Null-värden 1
4273 Null-värdet 1
4274 Numera 2
4275 Numeriska 1
4276 Nuova 1
4277 Nuts 1
4278 Nuvarande 1
4279 Nya 8
4280 Nyckeln 1
4281 Nyexploaterade 1
4282 Nyheterna 1
4283 Nyligen 2
4284 Nyss 1
4285 Nytt 2
4286 Nyttan 2
4287 Nyttofordon 1
4288 Nz 2
4289 Nämnda 1
4290 När 342
4291 Nära 1
4292 Näringslivet 1
4293 Närmare 2
4294 Nästa 84
4295 Nästan 3
4296 Nå 3
4297 Någon 17
4298 Någonstans 1
4299 Någonting 4
4300 Något 12
4301 Några 19
4302 Nåja 3
4303 Nån 1
4304 Nåväl 3
4305 Nödvändigheten 1
4306 Nödvändigt 1
4307 Núñez 1
4308 O 1
4309 OAS 1
4310 OAU 2
4311 OAVHÄNGIGHETEN 1
4312 OCH 2
4313 OCHA 1
4314 OECD 2
4315 OECD-länderna 1
4316 OFSR 1
4317 OFÖRBÄTTRAD 1
4318 OK 1
4319 OLAF 20
4320 OLAF:s 1
4321 OLE 2
4322 OLFAF 1
4323 OM 2
4324 OMRÖSTNING 9
4325 OSSE 1
4326 OSSE-observatörer 1
4327 OSSE:s 1
4328 OTC-derivat 10
4329 OTC-derivaten 3
4330 OTC-instrument 6
4331 OTC-instrumenten 1
4332 OTC-investeringar 1
4333 Oanmälda 1
4334 Oansvarighet 1
4335 Oavsett 7
4336 Oavslutad 1
4337 Oberbayern 1
4338 Oberoende 4
4339 Obnova-programmen 1
4340 Obs 1
4341 Observera 1
4342 Och 293
4343 Också 12
4344 Odara 11
4345 Odaras 2
4346 Oddy 1
4347 Odysseus 1
4348 Offentliga 2
4349 Offentligheten 1
4350 Office 25
4351 Office-pivottabellkomponent 1
4352 Office-program 1
4353 Offret 1
4354 Ofta 4
4355 Oförfärat 1
4356 Oförmögna 1
4357 Oil 3
4358 Oil-programmet 1
4359 Ojala 1
4360 Ojeda 1
4361 Okej 1
4362 Oklahoma 1
4363 Olika 3
4364 Olivia 7
4365 Olivias 1
4366 Olivier 1
4367 Oljebälte 1
4368 Oljebältet 1
4369 Oljestället 1
4370 Oljetankern 1
4371 Oljeutsläppet 1
4372 Olle 4
4373 Olyckan 2
4374 Olyckligtvis 1
4375 Olympe 1
4376 Olympic 1
4377 Olympiska 1
4378 Om 403
4379 Omagh 1
4380 Omfattande 1
4381 Omfånget 1
4382 Omkring 1
4383 Omlastningar 1
4384 Omorganisation 1
4385 Omräknat 1
4386 Området 3
4387 Omröstningen 56
4388 Omstrukturering 2
4389 Omstruktureringen 1
4390 Omständigheterna 1
4391 Omyndiga 1
4392 Onabu 1
4393 Onesta 1
4394 Online 1
4395 Onödigt 1
4396 Oomen-Ruijten 1
4397 Oostlander 3
4398 Operators 1
4399 Opinionsnätverk 1
4400 Oppositorum 1
4401 Oraninvånarnas 1
4402 Ord 3
4403 Orden 2
4404 Order 1
4405 Orderdetaljer 1
4406 Orderingången 1
4407 Ordet 6
4408 Ordförande 9
4409 Ordföranden 3
4410 Ordförandeskap 1
4411 Ordförandeskapet 9
4412 Ordförandeskapets 2
4413 Organet 1
4414 Organisationen 2
4415 Organization 1
4416 Orienten 2
4417 Orkanen 2
4418 Orkney 1
4419 Ormen 1
4420 Oron 2
4421 Oroväckande 1
4422 Orsaken 6
4423 Orsakerna 1
4424 Ortega 4
4425 Orwell 2
4426 Osip 1
4427 Oslo 3
4428 Osloavtalen 2
4429 Osloprotokollet 1
4430 Osman 1
4431 Ospar 6
4432 Ospar-avtalen 1
4433 Ospar-konventionen 3
4434 Ospar-målen 2
4435 Ospar-målet 1
4436 Ospar-normen 1
4437 Ospar-värdet 1
4438 Ostindiska 1
4439 Osäkerhet 1
4440 Otaliga 1
4441 Otroligt 1
4442 Oturligt 1
4443 Otvivelaktigt 1
4444 Ouvrière 1
4445 Oxonian 1
4446 Oz 3
4447 PATH 1
4448 PNV 1
4449 PPE 5
4450 PPE-DE 6
4451 PPE-DE- 2
4452 PPE-DE-gruppen 3
4453 PPE-DE-gruppens 2
4454 PPE-DE-ledamöter 1
4455 PPE-gruppen 4
4456 PPE-gruppens 1
4457 PR-effekt 1
4458 PR-experter 1
4459 PR-firmor 1
4460 PSE 2
4461 PSE-gruppen 5
4462 PSE-gruppens 3
4463 PT 27
4464 PVC 3
4465 PVC-leksaker 1
4466 Pack 3
4467 Package 1
4468 Packs 2
4469 Padanien 2
4470 Paddington 2
4471 Page 2
4472 Pakistan 4
4473 Pakistans 1
4474 Palacio 18
4475 Palacios 2
4476 Palermo 1
4477 Palestina 10
4478 Palestina-Israel 1
4479 Palestinaflyktingarnas 1
4480 Palestinafrågan 1
4481 Palestinas 2
4482 Palestinierna 1
4483 Panama 1
4484 Panza 1
4485 Paolo 1
4486 Papandreou 1
4487 Papayannakis 3
4488 Papoutsis 1
4489 Pappa 2
4490 Paracelsus 1
4491 Paradoxalt 2
4492 Paragrafrytteriet 1
4493 Parallella 1
4494 Parallellt 2
4495 Paris 6
4496 Parisfördragen 1
4497 Parisprotokollet 1
4498 Park 3
4499 Parken 1
4500 Parker 1
4501 Parlament 2
4502 Parlamentet 95
4503 Parlamentets 8
4504 Parlamentsledamöterna 1
4505 Parlamentsledamöternas 1
4506 Parlement 1
4507 Partido 1
4508 Partnerskap 1
4509 Partnerskapet 1
4510 Partnerskapets 1
4511 Pas 1
4512 Passagerarna 1
4513 Patricia 1
4514 Patten 55
4515 Pattens 8
4516 Paul 9
4517 Paul-Marie 1
4518 Pays 1
4519 Pays-de-Loire 1
4520 Peake 2
4521 Pecunia 1
4522 Peijs 2
4523 Peking 2
4524 Pekingdeklarationen 1
4525 Pekingkonferensen 1
4526 Pen 1
4527 Pensioner 1
4528 Pensionsfonder 1
4529 Pensionärerna 1
4530 Pensionärspartiet 3
4531 Pentagon 1
4532 Percy 4
4533 Peres 1
4534 Perfomance 1
4535 Person 1
4536 Personalsystemet 1
4537 Personer 1
4538 Personligen 8
4539 Peter 12
4540 Peters 2
4541 Petersberg 2
4542 Petersberguppgifter 1
4543 Petersberguppgifterna 3
4544 Petersen 1
4545 Petroleum 1
4546 Pettigrew 5
4547 Pettigrews 2
4548 Petunia 11
4549 Petunias 4
4550 Phare 6
4551 Phare- 1
4552 Phare-programmen 1
4553 Phare-programmet 2
4554 Philippe 1
4555 Philoxenia-programmet 2
4556 Phonograms 1
4557 Piecyk 4
4558 Pietrasanta 1
4559 Pietro 9
4560 Pietro-betänkandet 1
4561 Pietros 4
4562 Pinochet 10
4563 Pinochet-Ugarte 1
4564 Pintassilgobetänkandet 1
4565 Piqué 1
4566 Pirker 1
4567 PivotChart-vyn 2
4568 PivotTable- 2
4569 PivotTable-vyn 1
4570 Pivotabellvyns 1
4571 Pivotdiagramvy 1
4572 Pivottabeller 2
4573 Pivottabellista 1
4574 Pivottabellvy 1
4575 Pjoska 1
4576 Places 1
4577 Plaid 1
4578 Planeringskommittén 1
4579 Planerna 1
4580 Plantation 1
4581 Plantin 1
4582 Plast- 1
4583 Plastindustrin 1
4584 Platon 1
4585 Platons 1
4586 Plenarsessionens 1
4587 Plooij-van 3
4588 Plumb 1
4589 Plumb-Delors-avtalet 1
4590 Pläderingen 1
4591 Plötsligt 4
4592 Poettering 11
4593 Poetterings 1
4594 Pohjamo 1
4595 Pojkaktig 1
4596 Pojkarna 1
4597 Pojken 4
4598 Polen 7
4599 Polens 1
4600 Polisen 2
4601 Poliser 1
4602 Polisstyrkan 1
4603 Political 1
4604 Politik 1
4605 Politiken 3
4606 Politikens 1
4607 Polje 1
4608 Pollution 3
4609 Polo 1
4610 Pomés 1
4611 Ponnambalam 1
4612 Poos 4
4613 Popo 1
4614 Popular 1
4615 Port 3
4616 Portugal 36
4617 Portugals 7
4618 Portuguesa 1
4619 Positiv 1
4620 Posselt 5
4621 Post 2
4622 Post-Europa 1
4623 Posten 4
4624 Postföretaget 1
4625 Postkontoren 1
4626 Postkontorets 1
4627 Postmarknaden 1
4628 Posts 1
4629 Postsektorn 2
4630 Posttjänsten 5
4631 Posttjänster 1
4632 Posttjänsterna 5
4633 Postverken 1
4634 Potentiella 1
4635 Potsdam 1
4636 Pottaskan 1
4637 Potter 4
4638 Poul 1
4639 Poulenc 1
4640 Power 4
4641 Prag 1
4642 Praktiskt 1
4643 Precis 18
4644 Premiärminister 1
4645 Premiärministrar 1
4646 Premiärministrarna 1
4647 Presentationen 1
4648 President 2
4649 Pressfrihet 2
4650 Presumtivt 1
4651 Preussag 1
4652 Principen 6
4653 Principförklaringar 1
4654 Prioriteringen 1
4655 Privatdetektiven 1
4656 Privatisering 1
4657 Privet 5
4658 Problem 2
4659 Problemen 3
4660 Problemet 19
4661 Procacci 2
4662 Procaccis 1
4663 Procentsatserna 1
4664 Processen 7
4665 Processer 1
4666 Processerna 1
4667 Prodi 103
4668 Prodi-dokument 1
4669 Prodi-kommissionen 1
4670 Prodikommissionen 1
4671 Prodis 26
4672 Producenten 1
4673 Producenternas 1
4674 Produkter 1
4675 Programmappen 1
4676 Programmen 3
4677 Programmet 8
4678 Projekt 1
4679 Projekten 2
4680 Projektet 1
4681 Prokollet 1
4682 Pronk 3
4683 Propaganda 1
4684 Property 2
4685 Protection 2
4686 Protocol 1
4687 Protokoll 1
4688 Protokollen 1
4689 Protokollet 14
4690 Provan 2
4691 Provans 1
4692 Príncipes 1
4693 Pröva 1
4694 Puddingen 1
4695 Puerta 2
4696 Punkt 4
4697 Purvis 4
4698 Putin 2
4699 Putins 1
4700 Pyrenéerna 1
4701 PÅ 1
4702 På 173
4703 Påståendet 1
4704 Pétain 1
4705 Pöbelvälde 1
4706 QE2 2
4707 QE2:s 1
4708 Quebec 1
4709 Quecedo 3
4710 Queiro 1
4711 Queiró 1
4712 Quentin 1
4713 Quijote 9
4714 Quinn 117
4715 Quinns 3
4716 Quousque 1
4717 RC 1
4718 REP 2
4719 REVOKE 1
4720 RINA 3
4721 ROWS 1
4722 RSPB 1
4723 Ra-Ra 1
4724 Rabin 1
4725 Rabingruppen 1
4726 Racan 1
4727 Rachidi 1
4728 Rack 2
4729 Radio 4
4730 Radwan 4
4731 Rafael 4
4732 Rambeslutet 1
4733 Rambouillet 1
4734 Ramdirektivet 2
4735 Ramen 1
4736 Ramlah 1
4737 Ramprogrammet 1
4738 Ramvillkoren 2
4739 Randzio-Plath 4
4740 Randzio-Plaths 1
4741 Raninsy 1
4742 Rapkay 8
4743 Rapkaybetänkandet 1
4744 Rapkays 2
4745 Rapporten 4
4746 Ras 7
4747 Raschhofer 1
4748 Rasismen 1
4749 Rasistiska 2
4750 Ratificeringen 1
4751 Rato 1
4752 Rauf 2
4753 Ravenna 1
4754 Rayburnspis 1
4755 Raymond 1
4756 Reactor 1
4757 Reading 1
4758 Reaktionen 1
4759 Real 1
4760 Rebecca 6
4761 Rechar-programmet 1
4762 Redan 12
4763 Redarna 1
4764 Rederiet 1
4765 Reding 7
4766 Redings 2
4767 Redvers 1
4768 RefLibPaths-nyckel 2
4769 Referenser 2
4770 Reformen 6
4771 Reformering 1
4772 Reformeringen 1
4773 Reformerna 1
4774 Reformprocessen 2
4775 Regensburg 1
4776 Regeringarna 1
4777 Regeringen 6
4778 Regeringsförhandlingar 1
4779 Regeringskonferensen 2
4780 Regeringskonferensens 1
4781 Reginald 2
4782 Regionala 1
4783 Regionalpolitiken 1
4784 Regionen 2
4785 Regioner 1
4786 Regionerna 1
4787 Regionkommittén 2
4788 Regis 1
4789 Regler 2
4790 Regleringen 1
4791 Reglerna 1
4792 Reith 1
4793 Rekommendation 1
4794 Rektorn 1
4795 Relevant 1
4796 Religionen 1
4797 Remington 1
4798 Remora 1
4799 Rengie 2
4800 Rengies 1
4801 Rent 2
4802 Report 1
4803 ReportML 5
4804 ReportML-filen 1
4805 ReportML-format 1
4806 Representantgrupperna 1
4807 Republikaner 1
4808 Republiken 12
4809 Reserves 1
4810 Resolution 1
4811 Resolutionen 1
4812 Resolutionens 1
4813 Resolutioner 1
4814 Resolutionsförslag 4
4815 Resolutionsförslaget 1
4816 Resource 1
4817 Restaurant 1
4818 Resten 2
4819 Resterande 1
4820 Resterna 2
4821 Restore 1
4822 Resultat 2
4823 Resultaten 4
4824 Resultatet 10
4825 Resurser 1
4826 Retroaktiv 1
4827 Revideringen 1
4828 Revisionsrätten 5
4829 Rezala 2
4830 Rhen 1
4831 Rhendalen 1
4832 Rhenguld 2
4833 Rhenlandets 1
4834 Rhino 5
4835 Rhodesia 4
4836 Rhodesierna 1
4837 Rhone-Poulenc 1
4838 Rhône-Alpes 1
4839 Rialto 1
4840 Ricardo 1
4841 Richard 1
4842 Richterskalan 2
4843 Ries 1
4844 Rights 2
4845 Riis-Jørgensen 2
4846 Rika 1
4847 Riktlinjer 1
4848 Riktlinjerna 3
4849 Ringen 1
4850 Ringholm 2
4851 Rio 4
4852 Rio- 1
4853 Rio-konferensen 1
4854 Rioförklaringen 1
4855 Risken 3
4856 Ritt 1
4857 Riverside 5
4858 Road 2
4859 Robert 2
4860 Robertson 1
4861 Rocard 1
4862 Rocards 1
4863 Rode 1
4864 Roissys 1
4865 Rojos 1
4866 Roland 2
4867 Rollen 2
4868 Roly 7
4869 Rom 8
4870 Rom- 1
4871 Romano 10
4872 Romfördraget 3
4873 Romfördragets 1
4874 Romkonferensen 1
4875 Romkonventionerna 1
4876 Román 2
4877 Ron 32
4878 Ronald's 1
4879 Rons 8
4880 Roo 1
4881 Room 1
4882 Roosevelt 1
4883 Ropet 1
4884 Rosenberg 1
4885 Ross-on-Wye 1
4886 Roth-Behrendt 10
4887 Roth-Behrendts 1
4888 Rothe 2
4889 Rotterdam 3
4890 Round 2
4891 Roure 1
4892 Rover 2
4893 Royal 2
4894 Rugby 1
4895 Rugovas 1
4896 Ruhren 1
4897 Ruiz 1
4898 Rummet 2
4899 Rumänerna 1
4900 Rumänien 18
4901 Runt 3
4902 Rush 1
4903 Rusjailo 1
4904 Rwanda 1
4905 Ryska 1
4906 Ryssarna 2
4907 Ryssland 19
4908 Rysslands 7
4909 Ryttare 1
4910 Räcker 1
4911 Rädda 1
4912 Räkna 1
4913 Rätten 1
4914 Rättsstaten 1
4915 Rättssäkerheten 1
4916 Rättstillämpningen 1
4917 Rättvisa 2
4918 Råder 1
4919 Rådet 35
4920 Rådets 17
4921 Rådsmötet 1
4922 Rådsordföranden 1
4923 Rådsordförandeskapet 1
4924 Réunion 3
4925 Röda 2
4926 Rörande 3
4927 Rösta 1
4928 Rösterna 1
4929 Röstförklaringar 1
4930 Röstförklaringar- 1
4931 Rött 1
4932 Rübig 2
4933 Rübigs 1
4934 SA 3
4935 SA-kontot 1
4936 SAP 1
4937 SCRS 1
4938 SCRS-undersökningen 1
4939 SEK 1
4940 SEK(1998 3
4941 SEK(1999)1279 2
4942 SEK(99)0066 1
4943 SELECT 1
4944 SEM-2000 1
4945 SMAKAR 1
4946 SN 1
4947 SOLAS 1
4948 SPÖ 3
4949 SQL 21
4950 SQL-fråga 1
4951 SQL-frågeläge 11
4952 SQL-frågelägen 5
4953 SQL-frågelägena 1
4954 SQL-frågeläget 1
4955 SQL-frågor 1
4956 SQL-specifikationen 1
4957 SQL-syntax 1
4958 SQL-syntaxen 1
4959 SQL-uttryck 2
4960 SQL-uttrycken 1
4961 SS 1
4962 STOA 1
4963 SUD 1
4964 SUM-DISTINCT-Pris 1
4965 Sa 1
4966 Sacharovpriset 1
4967 Sadat 2
4968 Sadats 2
4969 Sages- 1
4970 Sagorna 1
4971 Sahara 4
4972 Sahel 1
4973 Saint-Exupérys 1
4974 Saint-Josse 1
4975 Sakellariou 1
4976 Sakellarious 1
4977 Saken 1
4978 Saker 2
4979 Salafranca 2
4980 Salafrancas 1
4981 Sam 4
4982 Samarbete 3
4983 Samarbetet 2
4984 Samarbetsavtalet 1
4985 Samband 1
4986 Sambandet 1
4987 Sambata 1
4988 Samhällena 1
4989 Samhället 2
4990 Samma 10
4991 Sammanfattningsvis 5
4992 Sammanflätningen 1
4993 Sammanhängande 1
4994 Sammanhållningen 1
4995 Sammanhållningsfonden 15
4996 Sammanhållningsfondens 1
4997 Sammansättningen 1
4998 Sammantaget 1
4999 Sammanträdena 1
5000 Sammanträdet 23
5001 Samordning 3
5002 Samordningen 1
5003 Samstämmighet 1
5004 Samstämmigheten 3
5005 Samtal 1
5006 Samtalen 1
5007 Samtidigt 43
5008 Samtliga 5
5009 San 2
5010 Sancho 1
5011 Sandbankar 1
5012 Sandbæk 1
5013 Sanningen 8
5014 Sanningens 1
5015 Sannolikt 1
5016 Santa 1
5017 Santer 3
5018 Santer-kommissionen 1
5019 Santer-kommissionens 1
5020 Santerkommissionens 1
5021 Santiago 1
5022 Santos 3
5023 Sapar 1
5024 Sapard 3
5025 Saramago 2
5026 Sardinernas 1
5027 Sarre-Lorraine-Luxemburg 1
5028 Saudiarabien 1
5029 Save 6
5030 Save- 1
5031 Save-programmet 2
5032 Savefloden 1
5033 Savimbi 1
5034 Savimbis 1
5035 Scabbers 1
5036 Scarborough 1
5037 Scenen 2
5038 Scharping 1
5039 Scheele 1
5040 Scheman 1
5041 Schengen 3
5042 Schengenavtalen 1
5043 Schengenavtalet 3
5044 Schengenkonventionen 1
5045 Schengenkonventionens 1
5046 Schengenområdet 1
5047 Schengenregelverket 1
5048 Schengenstat 1
5049 Scherers 1
5050 Schierhuber 1
5051 Schipol-flygplats 1
5052 Schleicher 3
5053 Schmid 1
5054 Schmidbetänkandet 1
5055 Schmidt 10
5056 Schmidtbetänkandet 1
5057 Schmidts 4
5058 Schori 2
5059 Schreyer 4
5060 Schroedter 10
5061 Schroedterbetänkandet 2
5062 Schroedters 6
5063 Schröder 1
5064 Schultz 2
5065 Schulz 7
5066 Schwaigerbetänkandet 1
5067 Schwarzwald 1
5068 Schweiz 3
5069 Schörling 1
5070 Schüssel 6
5071 Schüssels 1
5072 Sdot 1
5073 Se 7
5074 Sea 1
5075 Seattle 23
5076 Sebastian 1
5077 Secretary 1
5078 Sedan 72
5079 Sedvänjorna 1
5080 Segni 1
5081 Segura 1
5082 Seguro 1
5083 Seixas 6
5084 Sekelgammal 1
5085 Sektorn 1
5086 Sellafield 1
5087 Seminarier 1
5088 Sen 8
5089 Senare 6
5090 Senast 1
5091 Sens 1
5092 Sent 1
5093 Seppänen 1
5094 Ser 1
5095 Serbien 32
5096 Serbiens 4
5097 Seriösa 1
5098 Server 5
5099 Server-användaren 1
5100 Server-databas 1
5101 Server-databasen 5
5102 Servern 1
5103 Service 1
5104 Sett 1
5105 Sevilla 1
5106 Sex 3
5107 Sha'ananim 1
5108 Shahar 5
5109 Shaping 3
5110 Sharm 4
5111 Sharm-el-Sheik 1
5112 Sheets 1
5113 Shell 3
5114 Shepherdstown 3
5115 Shetland 1
5116 Shetlandsöarna 2
5117 Shimon 1
5118 Shinza 10
5119 Shinzas 1
5120 ShippedCity-fältet 1
5121 ShippedDate 1
5122 Shipping 2
5123 Shop 1
5124 Short 1
5125 Shropshire 1
5126 Sibirien 1
5127 Sicilien 1
5128 Siciliens 1
5129 Sid 1
5130 Side 1
5131 Sidor 1
5132 Siena 1
5133 Sierra 1
5134 Sifferuppgifterna 1
5135 Siffran 1
5136 Siffrorna 1
5137 Sihanouk 1
5138 Sikten 1
5139 Silver 4
5140 Simpson 1
5141 Sin 1
5142 Sinjavskij 2
5143 Sintra 8
5144 Sintraavtal 1
5145 Sintrafördraget 1
5146 Sion 1
5147 Sions 1
5148 Sir 2
5149 Siri 2
5150 Sist 2
5151 Sisyfosarbete 1
5152 Sisyfosklippa 1
5153 Sitting 1
5154 Situationen 15
5155 Sju 1
5156 Sjukdomen 3
5157 Sjukhusläkare 1
5158 Sjukvård 1
5159 Själv 5
5160 Själva 4
5161 Självfallet 1
5162 Självklart 6
5163 Sjätte 2
5164 Sjömäns 1
5165 Sjöstedt 7
5166 Sjötransporten 1
5167 Ska 3
5168 Skadestånd 1
5169 Skador 1
5170 Skadorna 1
5171 Skall 9
5172 Skapa 1
5173 Skapandet 3
5174 Skaror 1
5175 Skattedebiteringen 1
5176 Skatteharmonisering 1
5177 Skatterna 1
5178 Skeppet 1
5179 Sker 1
5180 Skickar 1
5181 Skillnaderna 3
5182 Skjulet 1
5183 Skogsvårdsmyndigheten 1
5184 Skopje 4
5185 Skotsk 1
5186 Skottland 25
5187 Skottlands 2
5188 Skrapie 1
5189 Skulden 1
5190 Skulle 26
5191 Skvallret 1
5192 Skydd 2
5193 Skyddet 4
5194 Skyddsåtgärderna 1
5195 Skyltar 1
5196 Skälen 1
5197 Skälet 6
5198 Slapphet 1
5199 Slovakien 1
5200 Slovenien 1
5201 Slut 1
5202 Sluta 1
5203 Slutligen 85
5204 Slutrapporten 1
5205 Slutresultatet 2
5206 Slutsatsen 3
5207 Slutsatserna 4
5208 Släpp 1
5209 Släppområden 3
5210 Släppområdena 1
5211 Slåss 1
5212 Smith 2
5213 Smiths 1
5214 Små 1
5215 Småföretagare 1
5216 Snabb 1
5217 Snarare 3
5218 Snart 3
5219 Snödrottningsspegel 1
5220 Soares 3
5221 Social 1
5222 Socialfonden 2
5223 Socialistgruppen 1
5224 Socialpolitik 1
5225 Socialpolitiken 2
5226 Socialpolitiska 1
5227 Society 1
5228 Soekarnopoetri 1
5229 Sokrates- 1
5230 Solana 52
5231 Solanas 4
5232 Solbes 6
5233 Soldat 1
5234 Soldater 1
5235 Solen 6
5236 Solidaritet 1
5237 Solidariteten 1
5238 Solsjenitsyns 1
5239 Som 183
5240 Somalia 1
5241 Somes 2
5242 Somliga 7
5243 Soppan 1
5244 Souchet 2
5245 Souladakis 2
5246 Southampton 2
5247 Souto 1
5248 Sovjetunionen 3
5249 Sovjetunionens 1
5250 Spanien 52
5251 Spaniens 4
5252 Spara 5
5253 Spararna 1
5254 Speciella 1
5255 Speciellt 1
5256 Specifika 2
5257 Spegelbilden 1
5258 Spelar 1
5259 Spencer 2
5260 Sperber 1
5261 Speroni 1
5262 Spindlarna 1
5263 Spinning 1
5264 Sport 1
5265 Spridda 1
5266 Språket 1
5267 Sputnikbaren 5
5268 Squeeze 1
5269 Sr 1
5270 Sri 3
5271 St 5
5272 Stabex- 1
5273 Stabiliserings- 1
5274 Stabiliteten 1
5275 Stabilitetspakten 3
5276 Stabilitetspaktens 1
5277 Stackars 5
5278 Staden 1
5279 Stadens 1
5280 Stadgan 3
5281 Stadsmiljöpolitiken 1
5282 Staes 1
5283 Stafford 1
5284 Stalins 1
5285 Standardinställningen 1
5286 Standardläge 1
5287 Standardläget 1
5288 Stanna 1
5289 Stapled 1
5290 Start- 1
5291 State 1
5292 Stater 1
5293 Staterna 6
5294 Staternas 1
5295 Station 1
5296 Stationerna 1
5297 Statistiken 1
5298 Statlig 1
5299 Statliga 2
5300 Statligt 1
5301 Statsbalen 1
5302 Statsmakten 1
5303 Steel 1
5304 Stegrennan 1
5305 Stegrennans 3
5306 Stegrennansstrandremsa 1
5307 Stella 6
5308 Stenar 1
5309 Stendhals 1
5310 Stenmarck 2
5311 Stenzel 8
5312 Stenzels 6
5313 Stephen 2
5314 Sterckx 5
5315 Stickordet 1
5316 Stilla 4
5317 Stillahavsområdet 2
5318 Stillman 54
5319 Stillmans 15
5320 Stjärnorna 1
5321 Stockholm 5
5322 Stoke-on-Trent 1
5323 Stolarna 1
5324 Stolen 1
5325 Stora 4
5326 Storbritannien 27
5327 Storbritanniens 2
5328 Storebror 1
5329 Storhertigdömet 1
5330 Storlek 1
5331 Stormar 1
5332 Stormarna 1
5333 Stormen 1
5334 Storskalig 1
5335 Stort 1
5336 Straffrätten 1
5337 Straffrättslig 1
5338 Straffrättsliga 1
5339 Straffångar 1
5340 Strasbourg 26
5341 Strasbourgförklaringen 2
5342 Strasbourgs 1
5343 Strategidokumentet 1
5344 Strategiska 1
5345 Stravinskij 1
5346 Strax 1
5347 Street 3
5348 Stregrennan 1
5349 Stromboli 2
5350 Strukturellt 2
5351 Strukturfonderna 2
5352 Strukturfondernas 2
5353 Sträckor 1
5354 Sträng 1
5355 Strävan 1
5356 Strävar 1
5357 Strålande 1
5358 Strömmen 1
5359 Studenter 1
5360 Studies 1
5361 Style 2
5362 Stylesheet 3
5363 Styrkan 1
5364 Städerna 1
5365 Stämmer 2
5366 Stämningen 2
5367 Ständiga 1
5368 Stålsektorn 1
5369 Ståndpunkterna 1
5370 Står 1
5371 Stöd 5
5372 Stöden 1
5373 Stöder 2
5374 Stödpunkten 1
5375 Stödsystemet 1
5376 Större 2
5377 Största 2
5378 Suanzes-Carpegna 4
5379 Subsidiariteten 1
5380 Subventioner 2
5381 Suckande 1
5382 Sudan 3
5383 Sudre 2
5384 Suffolk 1
5385 Sui 1
5386 Suicide 1
5387 Suisse 1
5388 Summan 1
5389 Suominen 2
5390 Suveräniteten 1
5391 Svaret 5
5392 Svart 1
5393 Svarta 1
5394 Svartvändargränden 2
5395 Svend 1
5396 Svenska 2
5397 Svepeskålen 1
5398 Sverige 44
5399 Sveriges 3
5400 Svårigheten 3
5401 Svårigheterna 1
5402 Svårt 1
5403 Swaziland 2
5404 Swedes 1
5405 Swoboda 15
5406 Swobodabetänkandet 1
5407 Swobodas 7
5408 Syd 8
5409 Sydafrika 24
5410 Sydafrikaavtalen 1
5411 Sydafrikas 2
5412 Sydamerika 2
5413 Sydeuropa 3
5414 Sydkorea 1
5415 Sydney 1
5416 Sydostasien 3
5417 Sydosteuropa 1
5418 Sydösteuropa 2
5419 Syftet 20
5420 Synd 1
5421 Synnerligen 1
5422 Syrien 27
5423 Syriens 2
5424 Syrierna 2
5425 Sysminsystemet 1
5426 Sysselsättningen 4
5427 Sysselsättningspakten 1
5428 Sysselsättningsstrategin 1
5429 System 1
5430 System32 1
5431 Systemadministratör 1
5432 Systemen 1
5433 Systemmappen 1
5434 Sánchez 3
5435 São 2
5436 Säg 2
5437 Säger 1
5438 Säker 1
5439 Säkerhet 1
5440 Säkerheten 1
5441 Säkerhetsaspekten 1
5442 Säkerhetskoefficienten 1
5443 Säkerhetsrådgivare 1
5444 Säkerhetsåtgärderna 1
5445 Säkerligen 2
5446 Säkert 1
5447 Sämre 1
5448 Särskild 2
5449 Särskilda 1
5450 Särskilt 12
5451 Säsongen 1
5452 Sättet 1
5453 Så 100
5454 Sådan 2
5455 Sådana 16
5456 Sådant 1
5457 Således 14
5458 Sålunda 3
5459 Såna 1
5460 Sången 1
5461 Sånt 2
5462 Såsom 9
5463 Såvitt 3
5464 Såväl 6
5465 Sète 1
5466 Söder 1
5467 Söderhavet 1
5468 Söderman 1
5469 Södermans 1
5470 Södern 1
5471 Sökvägarna 1
5472 Sörensen 1
5473 T-tack 1
5474 T.ex. 1
5475 T.o.m. 1
5476 TA 1
5477 TBT 3
5478 TDI-gruppen 3
5479 TILL 1
5480 TO 1
5481 TRIPS 1
5482 TRIPS-avtalen 2
5483 TSE 5
5484 TSE-risker 1
5485 TSE-sjukdomar 3
5486 TSQL 2
5487 TV 8
5488 TV-apparaten 1
5489 TV-apparater 1
5490 TV-bevakningen 1
5491 TV-bilder 1
5492 TV-bilderna 1
5493 TV-bolagen 1
5494 TV-kanal 4
5495 TV-kanalen 2
5496 TV-kanaler 3
5497 TV-program 2
5498 TV-programmen 1
5499 TV-skärmar 1
5500 TV-skärmen 1
5501 TV-sändare 1
5502 TV-team 1
5503 TV-tekniker 1
5504 TV-torn 1
5505 TV-utsändningar 1
5506 TV:n 1
5507 Ta 15
5508 Table 1
5509 Tacis 4
5510 Tacis- 1
5511 Tacis-programmet 2
5512 Tack 129
5513 Tadzjikistan 5
5514 Tag 1
5515 Taiwan 1
5516 Tajani 1
5517 Tajo-Segura- 1
5518 Tal 1
5519 Tala 2
5520 Talar 5
5521 Talaren 1
5522 Talisman 1
5523 Talmannen 24
5524 Tammerfors 33
5525 Tammerforsavtalen 1
5526 Tammerforsbeslutens 1
5527 Tang 1
5528 Tanganyika 1
5529 Tanio 1
5530 Tanken 5
5531 Tant 1
5532 Tanzania 2
5533 Tar 1
5534 Tarek 1
5535 Tas 1
5536 Tatu 1
5537 Tauerntunneln 1
5538 Taxis 1
5539 Tecken 1
5540 Teheran 1
5541 Tekniska 2
5542 Telefonen 1
5543 Telekommunikationsministeriet 1
5544 Telford 1
5545 Teresa 1
5546 Terror 1
5547 Terrorism 1
5548 Terroristerna 1
5549 Terrón 5
5550 Tesauro 1
5551 Texas 2
5552 Texten 3
5553 Thaci 1
5554 Thailand 1
5555 The 9
5556 Theato 12
5557 Theatobetänkandet 1
5558 Theatos 12
5559 Themsenmynningen 2
5560 Themsenvatten 1
5561 Theo 1
5562 Theonas 2
5563 Thermonuclear 1
5564 Thompson 1
5565 Thompsons 1
5566 Thors 3
5567 Thurber 1
5568 Thurn 1
5569 Thyssen 3
5570 Thyssens 2
5571 Tibet 22
5572 Tibet-frågan 1
5573 Tiden 2
5574 Tidigare 7
5575 Tidningsartiklarna 1
5576 Tidsfristen 2
5577 Tidsklyftan 1
5578 Tidvattnet 1
5579 Tiffanys 1
5580 Till 107
5581 Tillfälligheter 1
5582 Tillförlitliga 1
5583 Tillgänglig 1
5584 Tillgången 1
5585 Tillhörande 1
5586 Tillsammans 4
5587 Tillståndet 2
5588 Tillverkarna 2
5589 Tillverkningen 1
5590 Tillväxt 2
5591 Tillväxten 1
5592 Tillämpning 1
5593 Tillämpningen 2
5594 Tillåt 15
5595 TillåtBorttagning 1
5596 TillåtRedigering 1
5597 TillåtTillägg 1
5598 Tillåter 3
5599 Times 5
5600 Timor 4
5601 Timothy 6
5602 Tindi 2
5603 Tingesten 1
5604 Tio 2
5605 Tiotusentals 1
5606 Tisza 3
5607 Titanic 1
5608 Titley 2
5609 Titleys 1
5610 Titta 2
5611 Tja 2
5612 Tjeckien 2
5613 Tjeckiens 2
5614 Tjejen 2
5615 Tjernobyl 1
5616 Tjetjenien 15
5617 Tjetjenienpolitik 1
5618 Tjugo 2
5619 Tjuvars 1
5620 Tjänstekvaliteten 1
5621 Tjänsternas 1
5622 Tobin-skatt 1
5623 Today 1
5624 Toddyblom 1
5625 Todinskatten 1
5626 Tokyo 1
5627 Toledo 1
5628 Tolstoi 1
5629 Tom 1
5630 Tomma 2
5631 Tomé 2
5632 Tongivande 1
5633 Tonvikten 3
5634 Tool 1
5635 Tools 1
5636 Toppmötena 1
5637 Toppmötet 5
5638 Torrey 3
5639 Torry 1
5640 Torsdag 1
5641 Torv 1
5642 Torven 1
5643 Total 8
5644 Total-Elf 1
5645 Total-Fina 3
5646 TotalFina 1
5647 Totaler 1
5648 Tour 1
5649 Toyota 1
5650 Trade-Related 1
5651 Tradition 1
5652 Traditionen 1
5653 Traditionsmässigt 1
5654 Trafalgar 1
5655 Trafiken 1
5656 Trafiksäkerheten 1
5657 Transact-SQL-kommandon 1
5658 Transformation 3
5659 Transitional 1
5660 Transnationella 1
5661 Transport 1
5662 Transportsäkerheten 1
5663 Trastfältet 1
5664 Travel 1
5665 Tre 7
5666 Treaty 2
5667 Tredje 1
5668 Trentin 1
5669 Trepca 1
5670 Tretti 1
5671 Trettiotre 1
5672 Trevligt 1
5673 Trident 2
5674 Tridentbasen 1
5675 Trittin 1
5676 Tro 1
5677 Trojkan 1
5678 Trolla 1
5679 Trollkarlar 1
5680 Tror 13
5681 Trots 46
5682 Trovärdigheten 2
5683 Trycket 1
5684 Trygghetsfrågor 1
5685 Träd 1
5686 Trädgården 1
5687 Tsatsos 6
5688 Tulsa 1
5689 Tunisien 1
5690 Tupperware 1
5691 Tupperwarekvällar 1
5692 Turin 1
5693 Turism 3
5694 Turismen 8
5695 Turismens 1
5696 Turistpolitiken 1
5697 Turkiet 72
5698 Turkiets 15
5699 Turkmenistan 2
5700 Tusen 1
5701 Tusentals 1
5702 Tvillingarnas 1
5703 Tvärs 1
5704 Tvärt 2
5705 Tvärtom 13
5706 Två 18
5707 Tvåtusen 1
5708 Ty 16
5709 Tycker 3
5710 Tyckte 1
5711 Tydliga 1
5712 Tydligen 2
5713 Tydligt 1
5714 Tyskland 40
5715 Tysklands 2
5716 Tystnaden 1
5717 Tyvärr 36
5718 Tänk 13
5719 Tänker 2
5720 Tåget 3
5721 Tågkraschen 1
5722 U 4
5723 U-länderna 1
5724 U-ländernas 1
5725 UCITS 4
5726 UCITS-direktivet 1
5727 UCK 5
5728 UCK-ledaren 1
5729 UCK:s 2
5730 UCLAF 1
5731 UDB 2
5732 UEN 1
5733 UEN-gruppen 3
5734 UNCTAD 1
5735 UNEF 1
5736 UNHCR 1
5737 UNIFIL 1
5738 UNITA 2
5739 UNITA-flygplatserna 1
5740 UNITA:s 2
5741 UNMIK 6
5742 US-dollar 1
5743 USA 36
5744 USA:s 2
5745 USD 1
5746 Uganda 1
5747 Ugglan 1
5748 Ukraina 2
5749 Ulster 2
5750 Undantag 1
5751 Undantagen 1
5752 Undantaget 1
5753 Under 110
5754 Underbart 1
5755 Underformulär 2
5756 Underlaget 1
5757 Underpunkten 1
5758 Undersökningarna 1
5759 Undvik 1
5760 Unga 1
5761 Ungdoms- 1
5762 Ungefär 2
5763 Ungern 6
5764 Ungerns 1
5765 Unice 2
5766 Unicef 1
5767 Unilever 1
5768 Union 2
5769 Unionen 24
5770 Unionens 5
5771 United 1
5772 Universal 1
5773 Universum 1
5774 Uppassare 1
5775 Uppbyggnaden 1
5776 Uppdateringen 1
5777 Uppenbarligen 3
5778 Uppfylls 1
5779 Uppföljning 2
5780 Uppgiften 3
5781 Uppgifterna 1
5782 Uppgiftslämnare 1
5783 Uppgörelsen 1
5784 Upphovsmannarättigheter 1
5785 Upphovsrättsinnehavare 1
5786 Upplysningens 1
5787 Uppriktigt 2
5788 Upprättandet 2
5789 Uppsikt 1
5790 Ur 19
5791 Urba- 1
5792 Urban 27
5793 Urban-betänkandet 1
5794 Urban-dagordning 1
5795 Urban-initiativ 1
5796 Urban-initiativet 6
5797 Urban-initiativets 1
5798 Urban-program 1
5799 Urban-programmen 1
5800 Urban-programmet 12
5801 Urban-projekten 4
5802 Urban-utvecklingspolitik 1
5803 Urbans 1
5804 Urquiola 2
5805 Ursprungligen 1
5806 Ursprungsbefolkningen 2
5807 Ursprungstexten 1
5808 Ursula 2
5809 Ursäkta 7
5810 Uruguayrundan 2
5811 Urvalskriterierna 1
5812 Usted 1
5813 Ut 1
5814 Utan 20
5815 Utanför 3
5816 Utarbetandet 1
5817 Utarmningen 1
5818 Utbildning 1
5819 Utbildningen 1
5820 Utbildningsministeriet 1
5821 Utdelningen 1
5822 Utestående 1
5823 Utflödet 1
5824 Utformningen 3
5825 Utförande 1
5826 Utgiften 1
5827 Utgifterna 1
5828 Utifrån 5
5829 Utkastet 2
5830 Utmaningarna 1
5831 Utmaningen 3
5832 Utmattad 1
5833 Utmärkt 3
5834 Utnyttjandet 1
5835 Utnämning 1
5836 Utnämningen 1
5837 Utom 1
5838 Utomjordingar 1
5839 Utseende 1
5840 Utskottet 24
5841 Utskottets 1
5842 Utsläppet 1
5843 Uttalande 1
5844 Uttalandena 1
5845 Uttjänta 1
5846 Uttryck 1
5847 Uttrycket 1
5848 Utvecklandet 1
5849 Utvecklaren 1
5850 Utvecklingen 5
5851 Utvecklingsländer 1
5852 Utvecklingspartnerskapen 2
5853 Utvecklingssamarbetets 1
5854 Utvidgning 2
5855 Utvidgningen 5
5856 Utvidgningens 1
5857 Utvärdera 1
5858 Utöver 3
5859 Uzbekistan 2
5860 V 7
5861 V-ställda 1
5862 V. 1
5863 VBA 1
5864 VD 1
5865 VEU 5
5866 VI 2
5867 VIII 2
5868 Vaclav 6
5869 Vad 265
5870 Vadan 1
5871 Valdez 1
5872 Valdez-katastrofen 2
5873 Valen 1
5874 Valencias 1
5875 Valentins 1
5876 Valet 3
5877 Valette 1
5878 Valle 1
5879 Vallelersundi 4
5880 Vallonien 1
5881 Valverdes 1
5882 Van 15
5883 Vandamaffärerna 1
5884 Vanligen 1
5885 Vanligtvis 1
5886 Vanurå 1
5887 Vapen 1
5888 Var 28
5889 Vare 4
5890 Varela 4
5891 Varelsen 1
5892 Varenda 3
5893 Varför 55
5894 Varifrån 1
5895 Varje 41
5896 Varken 7
5897 Varning 1
5898 Varor 1
5899 Vart 3
5900 Vatanen 3
5901 Vatikanen 2
5902 Vatten 12
5903 Vattenbruket 1
5904 Vattenfrågan 1
5905 Vattenproblemet 1
5906 Vattnet 6
5907 Vautrin-beundrande 1
5908 Velzen 2
5909 Vem 25
5910 Vems 2
5911 Vendée 6
5912 Venetia 4
5913 Venezuela 2
5914 Venstres 2
5915 Ventimiglia 1
5916 Verheugen 8
5917 Verkligheten 2
5918 Verksamheten 2
5919 Verksamhetsområdet 1
5920 Verktyg 1
5921 Verktyg-menyn 1
5922 Vermeers 1
5923 Vernon 24
5924 Vernons 4
5925 Versailles 2
5926 Verts 4
5927 Verts-gruppens 1
5928 Vet 2
5929 Vetenskapen 1
5930 Vetenskapsmännen 2
5931 Veteranbilarnas 1
5932 Vetskapen 1
5933 Vi 1673
5934 Via 5
5935 Vice 1
5936 Viceconte 6
5937 Vicecontes 4
5938 Vichy-regeringens 1
5939 Vichyregimens 1
5940 Vid 63
5941 Vidal-Quadras 1
5942 Vidare 27
5943 Vietnams 1
5944 Vigo 1
5945 Vikten 1
5946 Viktiga 4
5947 Viktigast 3
5948 Vilagarcia 1
5949 Vild 1
5950 Vilda 2
5951 Viljan 1
5952 Vilka 39
5953 Vilken 17
5954 Vilket 7
5955 Vill 15
5956 Ville 2
5957 Villiers 5
5958 Villkoren 2
5959 Villkorliga 1
5960 Villkorsstyrd 1
5961 Vilse 1
5962 Vin 1
5963 Vinci 2
5964 Vinden 2
5965 Vinet 1
5966 Vinter 1
5967 Vintergatan 3
5968 Viout 1
5969 Vireaid 1
5970 Virginia 11
5971 Viruset 2
5972 Visa 4
5973 Vissa 34
5974 Visserligen 7
5975 Visst 11
5976 Visual 3
5977 Vit 1
5978 Vita 1
5979 Vitboken 3
5980 Vitheten 1
5981 Vitoria 2
5982 Vitorino 13
5983 Vitorinos 4
5984 Vivianne 1
5985 Vivien 6
5986 Vivienne 1
5987 Vlaams 1
5988 Vlaamsblok 1
5989 Vladimir 3
5990 Vodafone-Mannesmann 1
5991 Voinet 1
5992 Vojvodina 1
5993 Voldemort 5
5994 Voldemorts 2
5995 Volksunie 1
5996 Volkswagen 1
5997 Von 1
5998 Vore 1
5999 Vraket 1
6000 VÄNNER 1
6001 Vägen 3
6002 Vägkontroller 1
6003 Väldigt 1
6004 Välj 1
6005 Väljer 2
6006 Välkommen 1
6007 Välkomsthälsning 3
6008 Vänstern 1
6009 Vänsterns 1
6010 Vänta 1
6011 Väntade 1
6012 Väntar 1
6013 Värden 1
6014 Värderade 2
6015 Världen 2
6016 Världens 1
6017 Världsbanken 4
6018 Världsbankens 1
6019 Världshandelsorganisationen 8
6020 Världshandelsorganisationens 5
6021 Världshälsoorganisationen 1
6022 Världshälsoorganisationens 2
6023 Världsnaturfonden 3
6024 Världspostföreningens 1
6025 Världssamfundet 2
6026 Värmen 1
6027 Västafrika 1
6028 Västatlantens 1
6029 Västbanken 4
6030 Västeuropa 1
6031 Västeuropeiska 3
6032 Västfrika 1
6033 Västindien 5
6034 Västmakterna 1
6035 Västprovinsen 1
6036 Västra 1
6037 Västsahara 1
6038 Västtyskland 1
6039 Västtysklands 1
6040 Växthuseffekten 1
6041 Våld 1
6042 Våldet 2
6043 Vår 57
6044 Våra 19
6045 Vårt 19
6046 Véronique 1
6047 W3C 3
6048 WCT 1
6049 WHERE 1
6050 WHO 1
6051 WINNT 1
6052 WIPO 5
6053 WIPO-avtalen 5
6054 WIPO-avtalet 10
6055 WIPO-fördragen 1
6056 WIPO-församlingen 1
6057 WIPO-överläggningar 1
6058 WIPO:s 1
6059 WPPT 1
6060 WTO 12
6061 WTO-förenlig 1
6062 WTO-förhandlingarna 1
6063 WTO-systemet 1
6064 WTO:s 5
6065 WWF 1
6066 Waddenzee 1
6067 Waffen 1
6068 Waffen-SS:s 1
6069 Wagners 1
6070 Wahid 2
6071 Wales 18
6072 Wall 1
6073 Wallström 16
6074 Wallströms 2
6075 Walter 2
6076 Warszawa 1
6077 Warszawapaktens 1
6078 Warszawas 1
6079 Washington 5
6080 Washingtons 3
6081 Watch 2
6082 Waterfold 1
6083 Watergates 1
6084 Watts 1
6085 Weasley 30
6086 Weasleys 8
6087 Web 10
6088 Webbsidans 1
6089 Weiler 1
6090 Weimarrepublikens 1
6091 Wellington 1
6092 Wentz 19
6093 Wentz' 1
6094 West 3
6095 Westminster 1
6096 Where 1
6097 Wide 5
6098 Wiebenga 2
6099 Wieland 4
6100 Wien 4
6101 Wijkman 2
6102 Wijkmans 2
6103 Wilhelmshaven 1
6104 William 5
6105 Wilson 4
6106 Wilsons 1
6107 Wiltshire 1
6108 Windows 7
6109 Windows-registret 1
6110 Winwardöarna 2
6111 Witness 1
6112 Wogau 18
6113 Wogaubetänkandet 1
6114 Wogaus 3
6115 Wolfsonstiftelsen 1
6116 Women 1
6117 Word 1
6118 Work 1
6119 Work-romanerna 1
6120 World 9
6121 Wray 1
6122 Wulf-Mathies 5
6123 Wuori 1
6124 Wurtz 10
6125 Wye 1
6126 Wye-avtalen 1
6127 Wye-avtalet 1
6128 Wynn 1
6129 Wyre 1
6130 X 1
6131 XI 2
6132 XML 18
6133 XML- 4
6134 XML-aktiverade 1
6135 XML-baserade 2
6136 XML-baserat 1
6137 XML-data 6
6138 XML-datadokument 2
6139 XML-definierade 1
6140 XML-dokument 20
6141 XML-dokumentet 1
6142 XML-element 1
6143 XML-fil 5
6144 XML-filer 2
6145 XML-informationen 2
6146 XML-källan 1
6147 XML-liknande 1
6148 XML-märken 2
6149 XML-protokollet 1
6150 XML-relaterade 1
6151 XML-schemafil 2
6152 XML-schemastandarden 2
6153 XML-standardformat 1
6154 XML-syntax 1
6155 XML-syntaxen 1
6156 XP 5
6157 XP-licens 5
6158 XP-licenser 1
6159 XP-nätverkslicens 1
6160 XP-program 2
6161 XSD 4
6162 XSL 1
6163 XSL-fil 1
6164 XSL-formatmall 1
6165 XSL-formatmallar 1
6166 XSL-transformationsfil 1
6167 XSLT 6
6168 XX 1
6169 XXVII:e 1
6170 XXVIII:e 1
6171 Yam 1
6172 Yarmouth 1
6173 Yasir 1
6174 Yasser 1
6175 Yassir 1
6176 Yawlen 1
6177 Yawning 1
6178 Yeu 1
6179 Yom 1
6180 York 14
6181 Yorker 1
6182 Yorks 1
6183 Yorkshire 3
6184 You 1
6185 Youngblood 1
6186 Youth 1
6187 Youthstart 2
6188 Yr 1
6189 Yrkandet 1
6190 Yrkesutbildning 1
6191 Ytterligare 6
6192 Ytterst 2
6193 Yttersta 1
6194 Yttrandet 2
6195 Yttre 3
6196 Zaire 1
6197 Zakaria 1
6198 Zambia 3
6199 Zeeland 3
6200 Zeus 8
6201 Zimbabwe 1
6202 Zimeray 1
6203 Zimmerling 1
6204 Zion 1
6205 [ 6
6206 ] 7
6207 _ 1
6208 a 19
6209 abonnentförteckningen 1
6210 absolut 127
6211 absoluta 7
6212 absorberad 1
6213 absorberade 2
6214 abstrakt 3
6215 absurd 3
6216 absurda 2
6217 absurditet 1
6218 absurt 5
6219 acceleration 1
6220 accelerator 1
6221 accelererad 1
6222 accelererande 1
6223 accent 1
6224 accentuerar 1
6225 accentueras 2
6226 accentueringarna 1
6227 acceptabel 2
6228 acceptabelt 8
6229 acceptabla 1
6230 acceptans 6
6231 acceptansen 2
6232 acceptansnivån 1
6233 acceptera 60
6234 accepterad 1
6235 accepterade 5
6236 accepterande 3
6237 accepterandet 1
6238 accepterar 18
6239 accepteras 18
6240 accepterat 7
6241 accepterats 5
6242 accountability 1
6243 ach 1
6244 ackumulerat 1
6245 acquis 3
6246 acquisition 1
6247 action 1
6248 ad 5
6249 adderar 1
6250 additionalitet 3
6251 additionaliteten 1
6252 additionalitets- 1
6253 additionalitetsprincipen 7
6254 additionella 3
6255 additiva 1
6256 adekvat 6
6257 adekvata 2
6258 adelsskap 1
6259 adjektiv 2
6260 adjektivet 1
6261 adjö 1
6262 administration 8
6263 administrationen 7
6264 administrationer 1
6265 administrativ 6
6266 administrativa 29
6267 administrativt 9
6268 administratörer 1
6269 administratörsgruppen 1
6270 administrera 1
6271 administreras 1
6272 adriatiska 3
6273 advokat 4
6274 advokaten 1
6275 advokater 2
6276 affischer 1
6277 affär 8
6278 affären 2
6279 affärer 8
6280 affärsbeslut 1
6281 affärsföretag 1
6282 affärsgrenar 1
6283 affärshemligheter 1
6284 affärslivets 1
6285 affärsmannahänder 1
6286 affärsmän 1
6287 affärsmännens 1
6288 affärsmässig 1
6289 affärspaketverksamhet 1
6290 affärsresor 1
6291 affärsrisker 2
6292 affärsstrukturer 1
6293 affärsstrukturerna 1
6294 afrikaner 3
6295 afrikanerna 1
6296 afrikansk 1
6297 afrikanska 13
6298 afrikanskt 3
6299 aftonskolan 1
6300 age 1
6301 agenda 6
6302 agendan 3
6303 agent 4
6304 agenterna 1
6305 agera 56
6306 agerade 2
6307 agerande 42
6308 agerandet 2
6309 agerar 15
6310 agerat 6
6311 agg 1
6312 agglomerationscentra 1
6313 aggregat 1
6314 aggregaten 1
6315 aggression 3
6316 aggressioner 1
6317 aggressiv 1
6318 aggressiva 2
6319 agitation 1
6320 agrara 1
6321 agronomisk 1
6322 agroturismen 1
6323 aid 1
6324 aids 10
6325 aids-situationen 1
6326 aidsbekämpning 1
6327 aidsepidemi 1
6328 aidspatienter 2
6329 aidsrelaterad 1
6330 aidsrelaterade 1
6331 aidssiffrorna 1
6332 aidsviruset 2
6333 ajournering 2
6334 akademisk 1
6335 akademiska 1
6336 akt 18
6337 akta 3
6338 aktat 1
6339 akten 1
6340 aktens 1
6341 akter 2
6342 akterna 3
6343 akterut 1
6344 akteröver 1
6345 aktie 1
6346 aktiebolag 1
6347 aktiebolagen 1
6348 aktiebolaget 3
6349 aktiebörserna 1
6350 aktiefonder 2
6351 aktieindex 1
6352 aktieinnehav 1
6353 aktieinvesteringar 1
6354 aktiekurserna 1
6355 aktiemarknaden 2
6356 aktiemarknader 1
6357 aktier 3
6358 aktierna 2
6359 aktieägare 3
6360 aktieägarna 2
6361 aktieägarnas 2
6362 aktion 6
6363 aktionen 2
6364 aktioner 7
6365 aktionerna 3
6366 aktionsgrupper 3
6367 aktionsgrupperna 1
6368 aktionsradie 1
6369 aktiv 23
6370 aktiva 15
6371 aktivare 5
6372 aktivera 3
6373 aktiverad 1
6374 aktiverar 1
6375 aktiveras 4
6376 aktivering 1
6377 aktivism 1
6378 aktivistiska 1
6379 aktivitet 10
6380 aktiviteten 2
6381 aktiviteter 13
6382 aktiviteterna 4
6383 aktiviteters 1
6384 aktivitetsbaserad 1
6385 aktivitetsbaserade 1
6386 aktivt 30
6387 aktning 2
6388 aktningsbetygelse 1
6389 aktningsvärda 2
6390 aktris 1
6391 aktualisera 2
6392 aktualiseras 2
6393 aktualisering 2
6394 aktuell 9
6395 aktuella 71
6396 aktuellare 2
6397 aktuellt 8
6398 aktör 3
6399 aktören 2
6400 aktörer 27
6401 aktörerna 18
6402 aktörernas 3
6403 aktörers 2
6404 akut 6
6405 akuta 8
6406 akvarelltonade 1
6407 akvarium 1
6408 akvavit 3
6409 al-Sharas 1
6410 alarmerande 4
6411 alban 1
6412 albaner 7
6413 albanerna 1
6414 albansk 2
6415 albanska 13
6416 albansktalande 1
6417 aldrig 155
6418 alert 1
6419 alf 1
6420 alfabetet 2
6421 alfabetets 1
6422 alfabetiseringsnivå 1
6423 alfer 1
6424 algbekämpning 1
6425 alias 3
6426 aliasnamn 1
6427 alibi 2
6428 alienist 1
6429 alkemiskt 1
6430 alkemister 1
6431 alkohol 8
6432 alkoholbeskattning 1
6433 alkoholen 1
6434 alkoholens 1
6435 alkoholhalten 1
6436 alkoholhaltiga 7
6437 alkoholkonsumtion 1
6438 alkoholkonsumtionen 3
6439 alkoholmissbruk 1
6440 alkoholmonopol 1
6441 alkoholmonopolet 2
6442 alkoholpolitiken 2
6443 alkoholprodukter 4
6444 alkor 1
6445 all 119
6446 alla 1255
6447 allas 21
6448 alldaglig 1
6449 alldeles 95
6450 allegorisk 1
6451 allegoriska 1
6452 allehanda 4
6453 allena 1
6454 allenarådande 1
6455 allergiska 1
6456 allesammans 13
6457 allestädes 1
6458 alleuropeisk 1
6459 alleuropeiskt 2
6460 allians 5
6461 alliansen 23
6462 allianser 2
6463 alliansfria 1
6464 allierad 2
6465 allierade 3
6466 allihop 5
6467 allihopa 1
6468 allmosor 2
6469 allmän 53
6470 allmängiltiga 1
6471 allmängiltigt 1
6472 allmänhet 44
6473 allmänheten 47
6474 allmänhetens 15
6475 allmänintresse 1
6476 allmänna 134
6477 allmännas 1
6478 allmänne 1
6479 allmännyttig 2
6480 allmännyttiga 7
6481 allmänpolitisk 1
6482 allmänt 57
6483 allokeringar 1
6484 allomfattande 1
6485 allra 40
6486 alls 83
6487 allsidig 2
6488 allsidigt 2
6489 allsmäktighet 1
6490 allt 636
6491 allteftersom 7
6492 alltfler 3
6493 alltför 134
6494 alltid 222
6495 alltifrån 3
6496 alltihop 15
6497 allting 19
6498 alltjämt 7
6499 alltmer 13
6500 alltsammans 10
6501 alltsedan 4
6502 alltså 191
6503 allvar 36
6504 allvaret 3
6505 allvarlig 37
6506 allvarliga 82
6507 allvarligare 11
6508 allvarligaste 6
6509 allvarligt 65
6510 allvarsamt 1
6511 alpackajacka 1
6512 alster 1
6513 alt 1
6514 altare 1
6515 alternativ 28
6516 alternativa 7
6517 alternativen 2
6518 alternativet 3
6519 alternativt 1
6520 amatördiplomati 1
6521 ambassad 1
6522 ambassadör 3
6523 ambassadören 1
6524 ambassadörer 3
6525 ambition 17
6526 ambitionen 7
6527 ambitioner 25
6528 ambitionerna 1
6529 ambitionernas 2
6530 ambitiös 19
6531 ambitiösa 22
6532 ambitiösare 2
6533 ambitiöse 1
6534 ambitiöst 10
6535 ambulans 1
6536 ambulanser 1
6537 amerikan 2
6538 amerikanarna 1
6539 amerikanen 1
6540 amerikaner 1
6541 amerikanerna 18
6542 amerikansk 6
6543 amerikanska 54
6544 amerikanske 1
6545 amerikanskt 2
6546 amfiteatraliskt 1
6547 amiraler 1
6548 ammunition 1
6549 amp 2
6550 an 20
6551 ana 7
6552 anade 2
6553 analogt 1
6554 analys 40
6555 analysen 10
6556 analyser 4
6557 analysera 21
6558 analyserar 1
6559 analyseras 5
6560 analyserat 3
6561 analyserna 1
6562 analytiskt 2
6563 anamma 3
6564 anammande 1
6565 anammar 1
6566 anammat 4
6567 anammats 1
6568 anar 1
6569 anblick 1
6570 anblicken 3
6571 anbudsförfarande 1
6572 anbudsförfaranden 1
6573 anbudsförfarandet 2
6574 anbudsgivare 1
6575 anbudsgivningen 1
6576 anbudsinfordran 2
6577 and 9
6578 anda 24
6579 andades 2
6580 andaluser 2
6581 andalusier 3
6582 andalusierna 1
6583 andalusiska 1
6584 andan 10
6585 andar 1
6586 andas 4
6587 ande 1
6588 andedräkt 2
6589 andel 15
6590 andelar 4
6591 andelen 7
6592 andemening 2
6593 andemeningen 5
6594 andens 1
6595 andetag 2
6596 andfådd 1
6597 andhämtningens 1
6598 andlig 1
6599 andliga 3
6600 andlige 1
6601 andra 1122
6602 andrabehandling 1
6603 andrabehandlingsrekommendation 5
6604 andrabehandlingsrekommendationen 5
6605 andrahandsbehandlingsrekommendation 1
6606 andrakammare 1
6607 andras 7
6608 andre 4
6609 andres 1
6610 anekdoter 1
6611 anemi 1
6612 anfall 2
6613 anfallen 2
6614 anföra 4
6615 anförande 21
6616 anföranden 15
6617 anförandena 3
6618 anförandet 3
6619 anföras 1
6620 anförs 2
6621 anfört 2
6622 anförtro 1
6623 anförtros 3
6624 anförtrott 1
6625 anförtrotts 2
6626 angav 3
6627 angavs 2
6628 ange 30
6629 angelägen 14
6630 angelägenhet 11
6631 angelägenheten 3
6632 angelägenheter 11
6633 angelägenheterna 1
6634 angeläget 9
6635 angelägna 12
6636 angelägnare 1
6637 angenäm 3
6638 angenämt 1
6639 anger 19
6640 anges 31
6641 angetts 2
6642 angivandet 2
6643 angivare 2
6644 angivarna 1
6645 angivelse 1
6646 angiven 1
6647 angiveri 1
6648 angivit 4
6649 angivna 2
6650 angjorde 1
6651 anglosaxiska 1
6652 angolaner 1
6653 angolanska 10
6654 angrep 2
6655 angrepp 9
6656 angreppen 1
6657 angreppet 1
6658 angreppskrig 1
6659 angreppssätt 4
6660 angripa 13
6661 angripas 2
6662 angripen 2
6663 angriper 4
6664 angrips 1
6665 angränsande 5
6666 angående 72
6667 angår 6
6668 angör 1
6669 anhopningen 1
6670 anhängare 9
6671 anhängiggjort 1
6672 anhängiggöranden 1
6673 anhålla 2
6674 anhållnas 1
6675 anhållne 1
6676 anhöriga 2
6677 aning 17
6678 aningar 1
6679 aningen 2
6680 aningslösa 1
6681 ankar 3
6682 ankare 1
6683 ankaret 2
6684 ankarplats 1
6685 anklaga 1
6686 anklagad 1
6687 anklagade 4
6688 anklagades 2
6689 anklagas 4
6690 anklagelse 1
6691 anklagelsen 2
6692 anklagelser 6
6693 anklagelserna 6
6694 anklarna 1
6695 anknutna 1
6696 anknytning 4
6697 anknyts 1
6698 ankommer 1
6699 ankomst 2
6700 ankomsten 3
6701 ankrade 2
6702 anlag 1
6703 anlagd 2
6704 anlagda 1
6705 anlagt 2
6706 anlagts 1
6707 anledning 79
6708 anledningar 9
6709 anledningarna 2
6710 anledningen 52
6711 anletsdrag 1
6712 anlitat 1
6713 anlägga 1
6714 anlägger 2
6715 anläggning 6
6716 anläggningar 5
6717 anläggningarna 2
6718 anläggningarnas 1
6719 anläggningen 3
6720 anläggningsarbeten 1
6721 anläggs 1
6722 anlända 3
6723 anlände 4
6724 anländer 1
6725 anlänt 3
6726 anlöpa 1
6727 anlöper 5
6728 anmodade 3
6729 anmodan 1
6730 anmodar 1
6731 anmäla 4
6732 anmälan 4
6733 anmälda 2
6734 anmäler 1
6735 anmälning 1
6736 anmälningar 2
6737 anmälningsplikt 3
6738 anmälningsplikten 1
6739 anmälningsplikter 1
6740 anmälningssystemet 3
6741 anmäls 2
6742 anmält 3
6743 anmälts 1
6744 anmärkning 13
6745 anmärkningar 8
6746 anmärkningarna 2
6747 anmärkningen 1
6748 anmärkningsvärd 3
6749 anmärkningsvärda 4
6750 anmärkningsvärt 6
6751 anmärkte 1
6752 annalkande 2
6753 annan 168
6754 annans 1
6755 annanstans 7
6756 annars 31
6757 annat 278
6758 annonsera 1
6759 annorlunda 27
6760 annorstädes 4
6761 anomali 1
6762 anonym 2
6763 anonyma 2
6764 anonymitet 1
6765 anordna 3
6766 anordnade 5
6767 anordnas 2
6768 anordnats 1
6769 anordning 4
6770 anordningar 3
6771 anpassa 27
6772 anpassad 9
6773 anpassade 9
6774 anpassas 14
6775 anpassat 5
6776 anpassats 1
6777 anpassbarhet 1
6778 anpassning 15
6779 anpassningar 5
6780 anpassningarna 3
6781 anpassningen 6
6782 anpassningsbarhet 2
6783 anpassningsetappen 1
6784 anpassningsfasen 1
6785 anpassningsförmåga 4
6786 anpassningsproblem 1
6787 anropa 1
6788 anrätta 1
6789 ansade 1
6790 ansamlingen 1
6791 ansats 4
6792 ansatsen 2
6793 ansatser 5
6794 ansatserna 1
6795 anse 10
6796 ansedda 1
6797 anseende 10
6798 ansenlig 3
6799 ansenliga 1
6800 ansenligt 1
6801 anser 500
6802 anses 24
6803 ansett 7
6804 ansikte 41
6805 ansikten 11
6806 ansiktena 3
6807 ansiktet 12
6808 ansiktshuden 1
6809 ansiktslöse 1
6810 ansiktsuttryck 2
6811 ansjovis 4
6812 ansjovisbestånden 6
6813 ansjovisbeståndet 3
6814 ansjovisen 1
6815 ansjovisfiske 1
6816 ansjovisfisket 2
6817 ansjoviskvoten 1
6818 ansjoviskvoter 1
6819 anskaffat 1
6820 anskaffning 2
6821 anskrämliga 1
6822 anslag 26
6823 anslagen 20
6824 anslaget 6
6825 anslagits 1
6826 anslagna 2
6827 anslagsbeviljandet 1
6828 anslagsförbrukning 1
6829 anslagsfördelningen 1
6830 anslogs 1
6831 ansluta 30
6832 anslutande 1
6833 anslutas 2
6834 ansluter 18
6835 anslutit 5
6836 anslutits 1
6837 anslutna 3
6838 anslutning 39
6839 anslutningar 1
6840 anslutningen 19
6841 anslutningsfil 18
6842 anslutningsfilen 9
6843 anslutningsfilens 1
6844 anslutningsfiler 1
6845 anslutningsförfarandet 3
6846 anslutningsförhandlingarna 6
6847 anslutningsinformationen 5
6848 anslutningsländerna 1
6849 anslutningsmedel 1
6850 anslutningsprocess 1
6851 anslutningsprojektet 1
6852 anslutningsstrategin 1
6853 ansluts 2
6854 anslå 4
6855 anslår 2
6856 anslås 4
6857 anslöt 2
6858 anspelade 2
6859 anspelningar 1
6860 anspråk 14
6861 anspråksfulla 1
6862 anspråkslösa 2
6863 anspråkslösaste 1
6864 anspråkslöshet 1
6865 anstrykning 1
6866 anstränga 8
6867 ansträngda 1
6868 ansträngde 5
6869 anstränger 10
6870 ansträngning 9
6871 ansträngningar 75
6872 ansträngningarna 11
6873 ansträngs 1
6874 ansträngt 5
6875 anställa 8
6876 anställande 1
6877 anställbara 1
6878 anställbarhet 6
6879 anställbarheten 2
6880 anställd 3
6881 anställda 38
6882 anställdas 8
6883 anställer 1
6884 anställning 10
6885 anställningarna 2
6886 anställningsförhållanden 1
6887 anställningskontrakt 1
6888 anställningsmöjligheter 1
6889 anställningsvillkor 1
6890 anställt 1
6891 anställts 1
6892 anständig 5
6893 anständiga 6
6894 anständighet 3
6895 anständigt 3
6896 anstår 1
6897 ansvar 220
6898 ansvara 6
6899 ansvarar 13
6900 ansvaret 76
6901 ansvarig 39
6902 ansvariga 53
6903 ansvarige 3
6904 ansvarigt 6
6905 ansvarsavgränsning 1
6906 ansvarsbefrielse 1
6907 ansvarsbefrielsen 1
6908 ansvarsbördor 1
6909 ansvarsfrihet 34
6910 ansvarsfriheten 7
6911 ansvarsfrihetsrapport 1
6912 ansvarsfrågan 3
6913 ansvarsfrågorna 1
6914 ansvarsfull 3
6915 ansvarsfulla 6
6916 ansvarsfullt 11
6917 ansvarsfyllda 1
6918 ansvarsfördelning 2
6919 ansvarsfördelningen 3
6920 ansvarsförhållandena 1
6921 ansvarskultur 1
6922 ansvarskännande 2
6923 ansvarskänsla 3
6924 ansvarsområde 7
6925 ansvarsområden 3
6926 ansvarsområdena 1
6927 ansvarsområdet 1
6928 ansvarsordning 1
6929 ansvarsposter 4
6930 ansvarstagande 2
6931 ansvarstagandet 1
6932 ansvarstilldelning 1
6933 ansvarsuppgifter 1
6934 ansåg 19
6935 ansågs 6
6936 ansöka 2
6937 ansökan 12
6938 ansökande 2
6939 ansökarland 2
6940 ansökarländer 4
6941 ansökarländerna 12
6942 ansöker 2
6943 ansökningar 3
6944 ansökningsbestämmelser 1
6945 ansökt 2
6946 anta 59
6947 antagande 8
6948 antaganden 3
6949 antagandeprocessen 1
6950 antagandet 21
6951 antagen 3
6952 antagit 25
6953 antagits 20
6954 antagligen 10
6955 antagna 6
6956 antal 141
6957 antalet 67
6958 antar 29
6959 antas 27
6960 ante 5
6961 ante-systemet 1
6962 antecknade 2
6963 antecknat 1
6964 anteckningar 1
6965 anteckningsblock 1
6966 anteckningsbok 2
6967 anteckningsboken 2
6968 antenner 2
6969 anti-europeisk 1
6970 anti-europeiska 1
6971 anti-gemenskapliga 1
6972 anti-irländska 1
6973 anti-rasistiska 1
6974 antibedrägerilagstiftning 1
6975 antibiotika 7
6976 antibiotikaresistensens 1
6977 antibiotikum 1
6978 antidemokratiska 1
6979 antidiskrimineringslagar 1
6980 antieuropeiska 2
6981 antifascist 1
6982 antifascistiska 2
6983 antifolklig 1
6984 antika 3
6985 antikaffär 1
6986 antikens 1
6987 antikolonialism 1
6988 antikryptogam 2
6989 antimögelmedel 1
6990 antingen 26
6991 antipersonella 2
6992 antisemitisk 1
6993 antisemitiska 2
6994 antisemitism 3
6995 antisociala 1
6996 antiterroristoperation 1
6997 antites 1
6998 antitrustbestämmelserna 1
6999 antog 42
7000 antogs 23
7001 antropogenisk 1
7002 antropolog 1
7003 antyda 2
7004 antydan 3
7005 antydas 1
7006 antydde 4
7007 antyddes 1
7008 antyder 7
7009 antytt 1
7010 antågande 1
7011 anvisade 1
7012 anvisning 1
7013 anvisningar 2
7014 anvisningarna 2
7015 använd 3
7016 använda 147
7017 användande 4
7018 användandet 1
7019 användare 12
7020 användaren 5
7021 användarens 1
7022 användares 2
7023 användargränssnitt 1
7024 användargränssnittet 3
7025 användarkonto 1
7026 användarkrav 1
7027 användarkraven 1
7028 användarna 4
7029 användarnamn 1
7030 användarnas 3
7031 användas 66
7032 användbar 4
7033 användbara 4
7034 användbarhet 1
7035 användbart 7
7036 använde 16
7037 använder 71
7038 användes 9
7039 användning 47
7040 användningar 1
7041 användningarna 1
7042 användningen 33
7043 används 63
7044 använt 12
7045 använts 13
7046 apartheid 1
7047 apartheid-ordning 1
7048 apelsin 1
7049 apos 1
7050 apostel 1
7051 apostrof 1
7052 apotek 1
7053 apoteket 1
7054 apparat 1
7055 apparaten 1
7056 apparater 2
7057 apparaterna 1
7058 appell 1
7059 appellationsdomstolen 1
7060 applicerade 1
7061 applicerar 2
7062 appliceras 2
7063 applicerats 1
7064 applikationer 2
7065 applåder 15
7066 applådera 1
7067 applåderade 1
7068 applåderar 3
7069 april 21
7070 apropå 3
7071 aptit 1
7072 arab 1
7073 araber 1
7074 araberna 2
7075 arabernas 1
7076 arabisk 2
7077 arabisk-israeliska 1
7078 arabiska 11
7079 arabstat 1
7080 arabstater 1
7081 arabvärlden 2
7082 arbeta 117
7083 arbetad 1
7084 arbetade 12
7085 arbetande 5
7086 arbetar 69
7087 arbetare 10
7088 arbetaren 1
7089 arbetarens 1
7090 arbetarklassens 1
7091 arbetarna 4
7092 arbetarnas 2
7093 arbetarpartis 1
7094 arbetarstadsdelar 1
7095 arbetas 1
7096 arbetat 30
7097 arbete 274
7098 arbeten 17
7099 arbetena 2
7100 arbetet 81
7101 arbetets 2
7102 arbets- 3
7103 arbetsanda 1
7104 arbetsaspekter 1
7105 arbetsavtal 2
7106 arbetsbelastning 1
7107 arbetsbeskrivningar 1
7108 arbetsbörda 4
7109 arbetsbördan 1
7110 arbetsdokument 4
7111 arbetsdokumenten 1
7112 arbetsformer 2
7113 arbetsfrågorna 1
7114 arbetsfördelning 2
7115 arbetsförhållanden 2
7116 arbetsförmedlingar 1
7117 arbetsförmedlingen 1
7118 arbetsförmåga 1
7119 arbetsgivare 10
7120 arbetsgivaren 2
7121 arbetsgivarens 2
7122 arbetsgivarna 2
7123 arbetsgivarnas 3
7124 arbetsgivarorganisationen 1
7125 arbetsgivarparti 1
7126 arbetsgrupp 17
7127 arbetsgruppen 3
7128 arbetsgrupper 4
7129 arbetsinkomster 1
7130 arbetsinsats 3
7131 arbetsinsatser 2
7132 arbetsinsatserna 1
7133 arbetsintensiva 2
7134 arbetskontraktet 1
7135 arbetskraft 14
7136 arbetskraften 7
7137 arbetskraftens 1
7138 arbetskraftsintensiva 2
7139 arbetskraftsrörlighet 1
7140 arbetskultur 2
7141 arbetskvalitet 2
7142 arbetslagstiftning 1
7143 arbetsliv 4
7144 arbetslivet 9
7145 arbetslivets 1
7146 arbetslösa 21
7147 arbetslösas 2
7148 arbetslöshet 37
7149 arbetslösheten 66
7150 arbetslöshetens 3
7151 arbetslöshetsersättningen 1
7152 arbetslöshetsnivåer 1
7153 arbetslöshetspolitik 1
7154 arbetslöshetsproblemet 2
7155 arbetslöshetssiffrorna 3
7156 arbetslöshetsunderstöd 1
7157 arbetsmarknad 8
7158 arbetsmarknaden 38
7159 arbetsmarknadens 16
7160 arbetsmarknaderna 2
7161 arbetsmarknadsfrågor 1
7162 arbetsmarknadsförhållandena 1
7163 arbetsmarknadslagarna 1
7164 arbetsmarknadsministern 1
7165 arbetsmarknadsministrar 1
7166 arbetsmarknadsmyndigheter 1
7167 arbetsmarknadsorganisationerna 1
7168 arbetsmarknadsparternas 1
7169 arbetsmarknadspolitik 1
7170 arbetsmarknadspolitiken 4
7171 arbetsmarknadsproblem 1
7172 arbetsmarknadsrelationer 1
7173 arbetsmetod 2
7174 arbetsmetoden 2
7175 arbetsmetoder 4
7176 arbetsmetoderna 3
7177 arbetsmigration 1
7178 arbetsmiljö 1
7179 arbetsmotivation 1
7180 arbetsmängd 1
7181 arbetsmässiga 1
7182 arbetsmöjligheter 1
7183 arbetsnormer 3
7184 arbetsnormerna 1
7185 arbetsoduglig 1
7186 arbetsområdet 2
7187 arbetsordning 5
7188 arbetsordningen 25
7189 arbetsorganisation 2
7190 arbetsorganisationen 2
7191 arbetsorganiseringen 1
7192 arbetsperiod 1
7193 arbetsplan 1
7194 arbetsplanen 5
7195 arbetsplaner 1
7196 arbetsplats 1
7197 arbetsplatsen 3
7198 arbetsplatser 14
7199 arbetsplatserna 2
7200 arbetsplikt 1
7201 arbetspost 1
7202 arbetsprocessen 1
7203 arbetsprogram 13
7204 arbetsprogrammet 4
7205 arbetsrelationerna 1
7206 arbetsrum 1
7207 arbetsrutiner 1
7208 arbetsrätt 1
7209 arbetsrätten 1
7210 arbetsrättsliga 1
7211 arbetssammanträde 1
7212 arbetsskapande 1
7213 arbetsstyrka 2
7214 arbetsstyrkan 1
7215 arbetssystem 1
7216 arbetssätt 1
7217 arbetssättet 1
7218 arbetssökande 1
7219 arbetstagare 46
7220 arbetstagaren 5
7221 arbetstagarens 1
7222 arbetstagares 4
7223 arbetstagarna 22
7224 arbetstagarnas 11
7225 arbetstid 2
7226 arbetstiden 6
7227 arbetstidens 1
7228 arbetstider 2
7229 arbetstidsdirektivet 2
7230 arbetstidsförkortning 3
7231 arbetstidskriterierna 1
7232 arbetstidsordning 1
7233 arbetstidsreglerna 1
7234 arbetstidsutformning 1
7235 arbetstillfällen 95
7236 arbetstillfällena 4
7237 arbetstillstånd 5
7238 arbetstillståndet 1
7239 arbetsuppgifter 4
7240 arbetsverktyg 1
7241 arbetsvillkor 7
7242 arbetsvillkoren 4
7243 arbetsvärlden 1
7244 arbetsyta 2
7245 are 1
7246 arena 1
7247 arenan 1
7248 arg 1
7249 argent 1
7250 argument 28
7251 argumentation 1
7252 argumentationen 1
7253 argumentationskraft 1
7254 argumenten 5
7255 argumentera 3
7256 argumenterar 3
7257 argumentet 4
7258 aristokrat 1
7259 arkeolog 1
7260 arkeologiska 1
7261 arkitekter 1
7262 arkitektur 1
7263 arkiv 1
7264 arkiveras 1
7265 arkiveringsbricka 1
7266 arkivutrymmen 1
7267 arm 4
7268 armar 4
7269 armarna 2
7270 armarnas 1
7271 armbandsur 1
7272 armbågarna 2
7273 armbåge 1
7274 armbågen 1
7275 armen 4
7276 armenierna 2
7277 armeniska 1
7278 armlängds 1
7279 armod 2
7280 armé 8
7281 armén 4
7282 arméns 2
7283 arrangemang 7
7284 arrangemangen 4
7285 arrangemanget 1
7286 arrangera 3
7287 arrangerandet 1
7288 arrangerat 1
7289 arrest 1
7290 arresterad 2
7291 arresterades 6
7292 arresterats 1
7293 arresteringar 3
7294 arrogans 1
7295 arrogant 1
7296 arroganta 2
7297 arsenal 1
7298 art 13
7299 arte 1
7300 artefakt 1
7301 arten 2
7302 arter 9
7303 arterna 3
7304 artificiell 1
7305 artificiella 1
7306 artig 1
7307 artiga 3
7308 artighet 3
7309 artighetsgest 1
7310 artigt 2
7311 artikel 236
7312 artikeln 1
7313 artiklar 10
7314 artiklarna 11
7315 artikulerade 1
7316 artister 1
7317 arton 5
7318 artonhundratalet 1
7319 artonhundratalsstil 1
7320 artärer 1
7321 arv 13
7322 arven 1
7323 arvet 3
7324 arvode 1
7325 arvoden 1
7326 arvsynden 1
7327 as 1
7328 asfalten 1
7329 asfalterade 1
7330 asiatiska 1
7331 ask 1
7332 aska 2
7333 askar 1
7334 asken 1
7335 askenasernas 1
7336 asket 1
7337 askkoppar 1
7338 asocial 1
7339 aspekt 18
7340 aspekten 15
7341 aspekter 51
7342 aspekterna 10
7343 aspirera 1
7344 assegajer 1
7345 assimilering 1
7346 assistans 1
7347 assistent 2
7348 assistenter 2
7349 assistenterna 4
7350 assistentstadga 1
7351 assisterad 1
7352 assistito 1
7353 associerade 4
7354 associeras 1
7355 associering 1
7356 associeringsavtal 9
7357 associeringsavtalen 2
7358 associeringsavtalet 6
7359 associeringsförfarande 1
7360 associeringsprocessen 2
7361 asterisk 1
7362 asteroid 1
7363 asteroiden 1
7364 astma 1
7365 astronomen 1
7366 astronomer 1
7367 astronomiska 1
7368 asyl 10
7369 asyl- 2
7370 asylbeslut 1
7371 asylfrågan 1
7372 asylförfarande 2
7373 asylförfarandet 1
7374 asylpolitik 1
7375 asylrätt 4
7376 asylsökande 18
7377 asylsökandena 1
7378 asymmetrierna 1
7379 asymmetriska 1
7380 at 2
7381 ateister 1
7382 atlantalliansen 1
7383 atlantfart 1
7384 atlantkusten 1
7385 atmosfär 5
7386 atmosfärens 1
7387 atomenergimyndigheten 1
7388 atomenergiorganet 2
7389 atomforskningscentret 1
7390 atomkraften 1
7391 atomkraftverk 1
7392 att 19203
7393 attack 2
7394 attacken 1
7395 attacker 7
7396 attackerna 1
7397 attentat 3
7398 attentatet 1
7399 attesterats 1
7400 attityd 17
7401 attityder 3
7402 attityderna 1
7403 attraktionskraft 1
7404 attraktiv 2
7405 attraktiva 3
7406 attraktivt 2
7407 attribut 3
7408 attributen 1
7409 atypiska 1
7410 atypiskt 1
7411 auctoritas 1
7412 audio-visuella 1
7413 audiovisuella 1
7414 auditorium 1
7415 augusti 5
7416 auktionerna 1
7417 auktorisation 3
7418 auktoriserad 1
7419 auktoriserade 1
7420 auktoriseringar 1
7421 auktoritativ 1
7422 auktoritet 7
7423 auktoriteter 1
7424 autofilter 2
7425 autofiltrering 2
7426 autografera 1
7427 automatik 2
7428 automatisk 1
7429 automatiska 2
7430 automatiskt 21
7431 autonoma 2
7432 autonomi 3
7433 autonomin 1
7434 autopilot 1
7435 av 8714
7436 avancera 2
7437 avancerade 2
7438 avancerat 2
7439 avant 2
7440 avart 1
7441 avbetalning 1
7442 avbrott 4
7443 avbrottet 5
7444 avbruten 3
7445 avbrutits 2
7446 avbrutna 1
7447 avbryta 2
7448 avbryter 5
7449 avbryts 2
7450 avbröt 11
7451 avbröts 13
7452 avböjer 1
7453 avdela 4
7454 avdelar 1
7455 avdelning 12
7456 avdelningar 4
7457 avdelningarna 1
7458 avdelningen 2
7459 avdelnings- 1
7460 avdemokratiserar 1
7461 avec 2
7462 avenyn 1
7463 aversion 1
7464 aveuropeisering 1
7465 avfall 39
7466 avfallet 15
7467 avfallets 1
7468 avfalls- 1
7469 avfallsdirektiven 1
7470 avfallsfisk 1
7471 avfallshantering 2
7472 avfallshanteringen 2
7473 avfallshanteringens 1
7474 avfallshanteringsavgift 1
7475 avfallsinsamlaren 1
7476 avfallsmängd 1
7477 avfallsström 1
7478 avfallsströmmar 2
7479 avfallsströmmarna 1
7480 avfallssystem 1
7481 avfallsämnen 1
7482 avfolkas 1
7483 avfolkats 1
7484 avfolkning 3
7485 avfolkningsbygder 1
7486 avfolkningsvåg 1
7487 avfälliga 1
7488 avfärd 1
7489 avfärdad 1
7490 avfärdade 2
7491 avförd 1
7492 avfördes 1
7493 avförs 1
7494 avförts 1
7495 avgaser 1
7496 avgav 2
7497 avge 7
7498 avger 6
7499 avges 1
7500 avgett 1
7501 avgick 5
7502 avgift 4
7503 avgifter 9
7504 avgiftsutjämning 1
7505 avgivit 1
7506 avgivits 1
7507 avgjorde 3
7508 avgjort 4
7509 avgjorts 2
7510 avgnimningen 1
7511 avgrund 1
7512 avgränsa 2
7513 avgränsade 3
7514 avgränsar 1
7515 avgränsat 1
7516 avgå 2
7517 avgående 1
7518 avgång 6
7519 avgångsåtgärder 1
7520 avgår 1
7521 avgått 1
7522 avgör 5
7523 avgöra 19
7524 avgörande 114
7525 avgörandet 2
7526 avgöras 4
7527 avgörs 5
7528 avhandla 1
7529 avhandlas 2
7530 avhandlats 1
7531 avhjälpa 3
7532 avhjälpande 1
7533 avhjälpas 1
7534 avhjälps 1
7535 avhjälpts 2
7536 avhänder 1
7537 avhängig 2
7538 avhängigt 2
7539 avhålla 2
7540 avhållit 1
7541 avigsidor 1
7542 aviserade 3
7543 aviserar 2
7544 aviseras 1
7545 aviserat 2
7546 aviserats 2
7547 avisering 1
7548 avkall 2
7549 avkastning 5
7550 avkastningen 3
7551 avkastningsdjur 1
7552 avklarad 2
7553 avklarats 1
7554 avkrok 1
7555 avkrävas 2
7556 avkrävt 1
7557 avkunnar 2
7558 avlade 2
7559 avlagd 1
7560 avlagringar 1
7561 avlagt 1
7562 avlastning 1
7563 avledda 2
7564 avleder 1
7565 avlida 1
7566 avlivad 1
7567 avlivar 1
7568 avlivas 1
7569 avlivning 1
7570 avloppet 2
7571 avloppshål 1
7572 avloppsrör 1
7573 avlutat 1
7574 avlyssna 1
7575 avlyssnas 1
7576 avlyssning 11
7577 avlyssningen 4
7578 avlyssningssystemet 1
7579 avlägga 2
7580 avlägsen 5
7581 avlägset 6
7582 avlägsna 22
7583 avlägsnade 2
7584 avlägsnande 2
7585 avlägsnandet 2
7586 avlägsnas 1
7587 avlägsnat 1
7588 avlämnats 1
7589 avlöses 1
7590 avlösning 1
7591 avmagringskur 1
7592 avmattning 2
7593 avnjöt 1
7594 avocadokärnan 1
7595 avocat 2
7596 avoghet 1
7597 avogt 1
7598 avpassade 1
7599 avprickning 1
7600 avrapportering 1
7601 avreglera 4
7602 avreglerad 5
7603 avreglerade 2
7604 avreglerar 2
7605 avregleras 2
7606 avreglerat 2
7607 avreglering 39
7608 avregleringar 1
7609 avregleringen 44
7610 avregleringens 1
7611 avregleringsetapp 3
7612 avregleringsfas 1
7613 avregleringsområdet 1
7614 avregleringspolitiken 1
7615 avregleringsprocess 1
7616 avregleringsprocessen 1
7617 avregleringsscenarierna 1
7618 avregleringssteget 1
7619 avresan 1
7620 avrinningsområde 1
7621 avrinningsområden 1
7622 avrunda 1
7623 avrätta 1
7624 avrättades 1
7625 avrättat 1
7626 avråda 1
7627 avröjda 1
7628 avsaknad 5
7629 avsaknaden 14
7630 avsatsen 2
7631 avsatt 3
7632 avsatta 3
7633 avsattes 2
7634 avsatts 3
7635 avse 4
7636 avsedd 9
7637 avsedda 13
7638 avseende 70
7639 avseenden 19
7640 avseendena 1
7641 avseendet 42
7642 avser 63
7643 avses 9
7644 avsett 16
7645 avsevärd 6
7646 avsevärda 11
7647 avsevärt 15
7648 avsides 3
7649 avsikt 62
7650 avsikten 11
7651 avsikter 16
7652 avsikterna 3
7653 avsiktlig 2
7654 avsiktliga 3
7655 avsiktligt 4
7656 avsiktsförklaring 1
7657 avsiktsförklaringar 2
7658 avskaffa 24
7659 avskaffade 3
7660 avskaffades 2
7661 avskaffande 4
7662 avskaffandet 3
7663 avskaffar 4
7664 avskaffas 1
7665 avskaffat 1
7666 avskaffats 1
7667 avsked 2
7668 avskeda 2
7669 avskedande 1
7670 avskedar 1
7671 avskedat 1
7672 avskilda 1
7673 avskiljas 1
7674 avskriva 1
7675 avskriver 1
7676 avskrivning 1
7677 avskruvad 1
7678 avskräcka 3
7679 avskräckande 2
7680 avskräckning 1
7681 avskräcks 1
7682 avskrädeshög 1
7683 avskuren 1
7684 avsky 5
7685 avskydd 1
7686 avskydde 1
7687 avskyr 1
7688 avskytt 1
7689 avskyvärda 3
7690 avskyvärt 1
7691 avskärma 2
7692 avskärmar 1
7693 avskärmat 1
7694 avskärmning 1
7695 avslag 2
7696 avslitet 1
7697 avslog 6
7698 avslogs 3
7699 avsluta 37
7700 avslutad 71
7701 avslutade 12
7702 avslutades 12
7703 avslutande 5
7704 avslutandet 1
7705 avslutar 10
7706 avslutas 12
7707 avslutat 9
7708 avslutats 4
7709 avslutning 6
7710 avslutningen 2
7711 avslutningsvis 13
7712 avslängd 1
7713 avslå 3
7714 avslår 1
7715 avslås 2
7716 avslöja 2
7717 avslöjade 3
7718 avslöjades 1
7719 avslöjande 3
7720 avslöjanden 1
7721 avslöjar 9
7722 avslöjas 1
7723 avslöjat 1
7724 avsmak 4
7725 avsmalnande 1
7726 avsnitt 8
7727 avsnitten 2
7728 avsnittet 4
7729 avspegla 1
7730 avspeglar 6
7731 avspeglas 7
7732 avspänd 1
7733 avspända 1
7734 avspänning 1
7735 avspärrningar 1
7736 avstamp 1
7737 avstannat 1
7738 avsteg 1
7739 avstod 6
7740 avstänga 1
7741 avstängde 1
7742 avstängning 2
7743 avstå 16
7744 avståenden 1
7745 avstånd 17
7746 avstånden 2
7747 avståndet 10
7748 avståndstagande 3
7749 avstår 7
7750 avstått 8
7751 avsägande 1
7752 avsätta 6
7753 avsättas 1
7754 avsätter 1
7755 avsättningarna 1
7756 avsåg 6
7757 avtacklade 1
7758 avtal 127
7759 avtalade 3
7760 avtalas 1
7761 avtalat 3
7762 avtalats 4
7763 avtalen 22
7764 avtalens 1
7765 avtalet 70
7766 avtalets 7
7767 avtals 1
7768 avtalsförbindelser 1
7769 avtalsinnehållet 1
7770 avtalslösning 1
7771 avtalspart 1
7772 avtalsparterna 2
7773 avtalsslutande 1
7774 avtalstexten 1
7775 avtalstexterna 1
7776 avtalsvillkoren 2
7777 avtar 1
7778 avtecknade 4
7779 avtecknat 1
7780 avtog 1
7781 avtvinga 1
7782 avund 1
7783 avundades 1
7784 avundas 2
7785 avundsjuka 1
7786 avundsvärda 1
7787 avvakta 5
7788 avvaktan 6
7789 avvaktande 2
7790 avvaktar 3
7791 avveckla 6
7792 avvecklas 4
7793 avvecklat 2
7794 avvecklats 1
7795 avveckling 3
7796 avverkningsklara 1
7797 avvika 1
7798 avvikande 4
7799 avvikelse 1
7800 avvikelser 4
7801 avviker 3
7802 avvisa 9
7803 avvisade 3
7804 avvisades 1
7805 avvisande 1
7806 avvisandet 1
7807 avvisar 6
7808 avvisas 1
7809 avvisat 3
7810 avvisats 2
7811 avvisning 2
7812 avvägd 4
7813 avvägning 4
7814 avvägningar 1
7815 avvägningen 1
7816 avvägningsfall 1
7817 avvägs 1
7818 avvägt 1
7819 avvänja 1
7820 avväpnade 1
7821 avvärja 3
7822 avyttring 1
7823 axel 2
7824 axeln 4
7825 axelryckning 3
7826 axla 1
7827 axlar 4
7828 axlarna 10
7829 b 8
7830 baby 1
7831 babyn 1
7832 bacill 1
7833 back-position 1
7834 backa 1
7835 backade 4
7836 backen 2
7837 backshish-mentalitet 1
7838 bad 16
7839 bada 2
7840 badar 1
7841 badet 1
7842 badhytterna 1
7843 badkaret 1
7844 badrummet 5
7845 badvattnet 1
7846 badwill 1
7847 bagage 2
7848 bagaget 1
7849 bagatell 1
7850 bagatelliserar 1
7851 bagatellisering 1
7852 bain 1
7853 bak 5
7854 bakad 1
7855 bakat 1
7856 bakbundna 1
7857 bakdanta 1
7858 bakdörren 4
7859 baken 1
7860 bakficka 1
7861 bakfönstret 1
7862 bakgata 1
7863 bakgrund 71
7864 bakgrunden 14
7865 bakgrundsförslag 1
7866 bakgrundsnivå 1
7867 bakgrundsutsläpp 1
7868 bakgrundsvärdena 2
7869 bakgård 1
7870 bakgårdar 1
7871 bakhåll 1
7872 bakifrån 2
7873 bakning 1
7874 bakom 101
7875 bakomliggande 6
7876 bakre 1
7877 baksidestext 1
7878 bakslag 1
7879 bakslaget 1
7880 bakslugt 1
7881 baksätet 3
7882 baktalade 1
7883 baktanken 1
7884 bakvägen 1
7885 bakvägspolitik 1
7886 bakåt 6
7887 bakåtsträvande 2
7888 bakåtverkande 1
7889 balans 45
7890 balansen 14
7891 balanser 2
7892 balansera 3
7893 balanserad 15
7894 balanserade 6
7895 balanserande 1
7896 balanserar 2
7897 balanseras 1
7898 balanserat 8
7899 balansering 1
7900 balansräkningar 1
7901 balansövning 1
7902 baldakinförsedda 1
7903 balen 3
7904 balkan 1
7905 ballader 1
7906 ballast 1
7907 ballon 1
7908 baltiska 1
7909 bana 4
7910 banalisera 2
7911 banaliserar 1
7912 banaliseringen 1
7913 bananbåtarna 1
7914 bananerna 1
7915 bananrepubliker 1
7916 banar 1
7917 banat 1
7918 banbrytande 1
7919 band 17
7920 banden 3
7921 banderoll 2
7922 bandet 3
7923 banditer 1
7924 bank 4
7925 banka 1
7926 bankade 2
7927 banken 1
7928 bankens 1
7929 banker 4
7930 banketter 1
7931 bankförvaltningen 1
7932 bankgarantier 5
7933 bankirer 2
7934 bankkoncernerna 1
7935 bankkonton 2
7936 bankrutt 2
7937 banksekretessen 1
7938 banksystemet 1
7939 bannlysningen 1
7940 bannlysts 1
7941 banor 3
7942 banshee 1
7943 bantas 1
7944 bantning 1
7945 bantningen 1
7946 bantningskur 1
7947 bar 21
7948 bara 882
7949 baracker 1
7950 barbari 1
7951 barbariet 2
7952 barbariets 1
7953 barbariska 2
7954 barbariskt 1
7955 barberarna 1
7956 baren 2
7957 barens 1
7958 barerna 1
7959 barkborren 1
7960 barm 3
7961 barn 74
7962 barn- 1
7963 barnadödlighet 4
7964 barnadödligheten 1
7965 barnafödande 1
7966 barnbarn 1
7967 barnbedrägeri 1
7968 barndom 1
7969 barndomen 2
7970 barndödlighet 3
7971 barndödligheten 1
7972 barnen 11
7973 barnens 8
7974 barnet 3
7975 barnets 1
7976 barnhandel 1
7977 barnhälsoproblemet 1
7978 barnmorska 1
7979 barnomsorg 2
7980 barnpornografi 2
7981 barns 6
7982 barnsligaste 1
7983 barnungar 1
7984 baron 1
7985 barriärer 2
7986 bars 4
7987 barskt 1
7988 bart 1
7989 bartender 1
7990 bas 6
7991 basackompanjemanget 1
7992 basar 2
7993 base 1
7994 baseball 1
7995 baseballmössor 1
7996 baseballresultaten 1
7997 basen 4
7998 baser 1
7999 basera 2
8000 baserad 6
8001 baserade 6
8002 baserar 4
8003 baseras 14
8004 baserat 7
8005 basförsörjning 1
8006 basis 6
8007 bask 4
8008 baskisk 3
8009 baskiska 12
8010 baskiskt 1
8011 baskolumnens 1
8012 baskrar 1
8013 basnivå 1
8014 bastardhunden 1
8015 bastu 1
8016 basunstöt 3
8017 basvattenförbrukning 1
8018 baxa 1
8019 bayerska 1
8020 bayerskt 1
8021 bayrare 1
8022 be 63
8023 beakta 29
8024 beaktades 5
8025 beaktande 7
8026 beaktanden 1
8027 beaktandet 2
8028 beaktansvärt 1
8029 beaktar 13
8030 beaktas 29
8031 beaktat 8
8032 beaktats 7
8033 bearbeta 2
8034 bearbetade 1
8035 bearbetande 1
8036 bearbetas 1
8037 beblandade 1
8038 bebodd 1
8039 bebodda 2
8040 bebyggelse 1
8041 bebyggelsen 1
8042 bebådade 1
8043 bedra 3
8044 bedragare 1
8045 bedragares 1
8046 bedrar 2
8047 bedrevs 1
8048 bedrifter 2
8049 bedriva 15
8050 bedrivas 5
8051 bedriver 12
8052 bedrivit 3
8053 bedrivs 7
8054 bedrägeri 15
8055 bedrägeribekämpning 7
8056 bedrägeribekämpningen 1
8057 bedrägerier 15
8058 bedrägerierna 1
8059 bedrägeriet 2
8060 bedrägerikonventionen 1
8061 bedrägerimål 1
8062 bedräglig 1
8063 bedrövelser 1
8064 bedrövliga 1
8065 bedrövligt 2
8066 bedöma 29
8067 bedömas 8
8068 bedömda 1
8069 bedömde 1
8070 bedömdes 1
8071 bedömer 11
8072 bedömning 41
8073 bedömningar 4
8074 bedömningarna 2
8075 bedömningen 8
8076 bedöms 9
8077 bedömt 2
8078 beef 1
8079 befallningar 1
8080 befann 9
8081 befara 2
8082 befarar 5
8083 befatta 2
8084 befattar 1
8085 befattat 4
8086 befattning 3
8087 befattningar 4
8088 befattningarna 1
8089 befinna 9
8090 befinner 92
8091 befintlig 2
8092 befintliga 51
8093 befintligt 1
8094 befläckad 1
8095 befogad 3
8096 befogade 3
8097 befogat 4
8098 befogenhet 11
8099 befogenheter 45
8100 befogenheterna 2
8101 befogenhetsområden 1
8102 befolka 1
8103 befolkad 1
8104 befolkade 6
8105 befolkning 34
8106 befolkningar 4
8107 befolkningarna 10
8108 befolkningarnas 2
8109 befolkningen 87
8110 befolkningens 10
8111 befolknings 1
8112 befolkningsdelar 1
8113 befolkningsgrupper 10
8114 befolkningsgrupperna 4
8115 befolkningskoncentration 1
8116 befolkningslager 1
8117 befolkningslagren 1
8118 befolkningsmajoriteten 2
8119 befolkningsmajoritetens 1
8120 befolkningssammansättningen 1
8121 befolkningssiffra 2
8122 befolkningsspridning 1
8123 befolkningsstorlek 1
8124 befolkningsstorleken 1
8125 befolkningsstruktur 1
8126 befolkningstillväxt 1
8127 befolkningstäthet 1
8128 befolkningstätheten 1
8129 befolkningsunderlag 1
8130 befordrad 1
8131 befordran 8
8132 befordras 1
8133 befraktare 1
8134 befraktaren 4
8135 befraktarna 2
8136 befraktarnas 3
8137 befria 1
8138 befriad 2
8139 befriar 1
8140 befrias 5
8141 befriat 2
8142 befriats 1
8143 befrukta 1
8144 befrämjandet 1
8145 befrämjat 1
8146 befullmäktigade 1
8147 befunnit 3
8148 befunnits 1
8149 befäl 2
8150 befälet 2
8151 befälhavare 2
8152 befälhavaren 1
8153 befängda 2
8154 befängt 1
8155 befäst 1
8156 befästa 11
8157 befästande 1
8158 befäste 1
8159 befäster 3
8160 befästes 1
8161 begagnade 6
8162 begav 1
8163 bege 3
8164 begrava 1
8165 begravning 3
8166 begravningsplatser 1
8167 begrep 2
8168 begrepp 17
8169 begreppen 5
8170 begreppet 32
8171 begripa 2
8172 begriper 4
8173 begriplig 1
8174 begripligare 1
8175 begripligt 3
8176 begrunda 3
8177 begrundade 1
8178 begränsa 42
8179 begränsad 38
8180 begränsade 28
8181 begränsades 2
8182 begränsande 2
8183 begränsar 19
8184 begränsas 17
8185 begränsat 15
8186 begränsats 1
8187 begränsning 12
8188 begränsningar 20
8189 begränsningarna 6
8190 begränsningen 1
8191 begränsningsavtal 1
8192 begynnande 1
8193 begynnelsebokstaven 1
8194 begynnelsen 2
8195 begynte 1
8196 begär 42
8197 begära 21
8198 begäran 63
8199 begäran.)Beträffande 1
8200 begäras 3
8201 begärda 1
8202 begärde 12
8203 begärets 1
8204 begärs 8
8205 begärt 24
8206 begå 3
8207 begångna 1
8208 begår 3
8209 begås 6
8210 begått 5
8211 begåtts 3
8212 begåvad 1
8213 begåvning 1
8214 behag 1
8215 behagligt 1
8216 behandla 36
8217 behandlad 1
8218 behandlade 5
8219 behandlades 6
8220 behandlar 38
8221 behandlas 50
8222 behandlat 10
8223 behandlats 4
8224 behandling 36
8225 behandlingarna 1
8226 behandlingen 50
8227 behandlingens 1
8228 behandlingsanläggning 1
8229 behandlingsanläggningarna 1
8230 behandlingscentraler 1
8231 behov 86
8232 behoven 12
8233 behovet 97
8234 behäftat 1
8235 behärskade 1
8236 behåll 1
8237 behålla 34
8238 behållare 1
8239 behållas 1
8240 behåller 2
8241 behållit 1
8242 behållits 1
8243 behålls 3
8244 behöll 3
8245 behölls 1
8246 behörig 2
8247 behöriga 15
8248 behörige 1
8249 behörighet 16
8250 behörigheten 2
8251 behörigheter 4
8252 behörighetsnivå 1
8253 behörighetsområde 4
8254 behörighetsområden 1
8255 behörigt 1
8256 behöva 52
8257 behövande 1
8258 behövas 6
8259 behövde 12
8260 behövdes 3
8261 behöver 268
8262 behövliga 1
8263 behövs 113
8264 behövt 3
8265 behövts 1
8266 beivras 1
8267 bekant 11
8268 bekanta 4
8269 bekantgjorts 1
8270 beklaga 20
8271 beklagade 3
8272 beklagande 6
8273 beklaganden 3
8274 beklagansvärd 1
8275 beklagansvärda 2
8276 beklagansvärt 3
8277 beklagar 49
8278 beklagat 2
8279 beklaglig 2
8280 beklagliga 3
8281 beklagligt 17
8282 beklämmande 2
8283 bekom 1
8284 bekostat 1
8285 bekostnad 7
8286 bekräfta 39
8287 bekräftade 5
8288 bekräftades 3
8289 bekräftande 1
8290 bekräftar 17
8291 bekräftas 9
8292 bekräftat 7
8293 bekräftats 4
8294 bekräftelse 5
8295 bekräftelsen 2
8296 bekväm 2
8297 bekvämligheter 2
8298 bekvämlighetsflagg 23
8299 bekvämlighetsflaggade 5
8300 bekvämlighetsflaggades 1
8301 bekvämlighetsflaggen 1
8302 bekvämlighetsflaggningen 1
8303 bekvämt 3
8304 bekymmer 17
8305 bekymmersamma 1
8306 bekymmersamt 3
8307 bekymra 1
8308 bekymrad 9
8309 bekymrade 8
8310 bekymrande 1
8311 bekymrar 7
8312 bekymrat 2
8313 bekämpa 76
8314 bekämpade 2
8315 bekämpande 3
8316 bekämpandet 2
8317 bekämpar 6
8318 bekämpas 3
8319 bekämpats 1
8320 bekämpning 13
8321 bekämpningen 5
8322 bekämpningsmedel 1
8323 bekänna 1
8324 bekännelse 1
8325 bekännelser 1
8326 bekänner 1
8327 belagda 1
8328 belagt 1
8329 belasta 1
8330 belastande 1
8331 belastar 2
8332 belastas 2
8333 belastning 4
8334 belastningar 1
8335 belgisk 3
8336 belgiska 13
8337 belopp 15
8338 beloppen 3
8339 beloppet 6
8340 beloppets 1
8341 belysa 2
8342 belysas 1
8343 belyser 2
8344 belysning 2
8345 belyst 2
8346 beläget 2
8347 belägg 1
8348 beläggs 1
8349 belägna 7
8350 belåtenhet 2
8351 belåtet 3
8352 belåtna 1
8353 belönar 1
8354 belönas 2
8355 belöpte 1
8356 bemannade 1
8357 bemanningsbehovet 1
8358 bemyndigande 6
8359 bemyndigar 1
8360 bemärkelse 4
8361 bemärkelsen 4
8362 bemästra 1
8363 bemöda 5
8364 bemödanden 4
8365 bemödar 1
8366 bemöta 10
8367 bemötande 1
8368 bemötas 1
8369 bemöter 5
8370 bemöts 2
8371 bemötts 1
8372 ben 11
8373 bench-marking 1
8374 benchmark 1
8375 benchmarking 3
8376 benchmarking-system 1
8377 benchmarks 1
8378 benen 5
8379 benet 1
8380 benhård 1
8381 benhårda 1
8382 benhårt 1
8383 benig 1
8384 benmjöl 1
8385 bensin 2
8386 bensinpriset 1
8387 benstomme 2
8388 benägna 3
8389 benämning 1
8390 benämns 1
8391 benåda 1
8392 beordra 1
8393 beordrat 1
8394 beordrats 1
8395 ber 104
8396 bereda 2
8397 beredas 1
8398 beredd 46
8399 beredda 44
8400 bereder 1
8401 beredningen 1
8402 bereds 1
8403 beredskap 3
8404 beredskapen 1
8405 beredvilligt 1
8406 berett 8
8407 beretts 2
8408 berg 6
8409 berget 2
8410 bergs- 1
8411 bergskommunerna 1
8412 bergsområden 1
8413 bergssektorer 1
8414 bergssidan 1
8415 berika 7
8416 berikande 2
8417 berikar 3
8418 berikas 1
8419 berikat 1
8420 bero 1
8421 berodde 6
8422 beroende 64
8423 beroendeminskning 1
8424 beroendet 3
8425 beror 55
8426 berott 2
8427 berusa 1
8428 berusad 2
8429 berusat 1
8430 beryktad 1
8431 beryktade 1
8432 beräkna 4
8433 beräknade 3
8434 beräknades 1
8435 beräknar 2
8436 beräknas 6
8437 beräknat 2
8438 beräknats 1
8439 beräkning 2
8440 beräkningar 5
8441 beräkningarna 4
8442 beräkningen 8
8443 berätta 28
8444 berättade 22
8445 berättar 6
8446 berättare 1
8447 berättas 1
8448 berättat 5
8449 berättelse 4
8450 berättelsen 3
8451 berättelser 1
8452 berättelserna 1
8453 berättiga 1
8454 berättigad 10
8455 berättigade 18
8456 berättigande 6
8457 berättigar 3
8458 berättigas 2
8459 berättigat 13
8460 berömd 3
8461 berömda 6
8462 berömde 1
8463 berömma 5
8464 berömmande 1
8465 berömt 1
8466 berömvärd 1
8467 berömvärda 2
8468 berömvärt 2
8469 berör 43
8470 beröra 2
8471 beröras 4
8472 berörd 2
8473 berörda 62
8474 berörde 4
8475 berördes 2
8476 beröring 1
8477 beröringen 1
8478 beröringspunkter 1
8479 berörs 21
8480 berört 8
8481 berörts 3
8482 beröva 3
8483 berövar 1
8484 berövats 1
8485 besatta 2
8486 besatthet 1
8487 besegla 1
8488 besegrade 1
8489 besegrades 1
8490 besegrar 1
8491 besiktning 1
8492 besiktningar 1
8493 besiktningsinstrument 1
8494 besiktningsmyndigheterna 1
8495 besitter 5
8496 beskaffenhet 1
8497 beskatta 2
8498 beskattad 1
8499 beskattas 1
8500 beskattning 9
8501 beskattningen 2
8502 beskattningsfrågor 1
8503 beskattningskod 1
8504 besked 12
8505 beskjuta 1
8506 beskrev 5
8507 beskrevs 3
8508 beskriva 12
8509 beskrivande 2
8510 beskrivas 3
8511 beskriver 11
8512 beskrivet 2
8513 beskrivit 9
8514 beskrivits 2
8515 beskrivna 2
8516 beskrivning 12
8517 beskrivningar 1
8518 beskrivs 11
8519 beskydd 6
8520 beskydda 1
8521 beskylla 1
8522 beskyller 1
8523 beskyllningar 1
8524 beskylls 1
8525 beskyllts 1
8526 beskåda 1
8527 besköt 1
8528 beslag 1
8529 beslagta 1
8530 beslagtagna 1
8531 beslut 265
8532 besluta 27
8533 beslutade 22
8534 beslutades 5
8535 beslutande 3
8536 beslutandefrihet 1
8537 beslutandemakten 1
8538 beslutandeplanet 1
8539 beslutanderätt 2
8540 beslutar 13
8541 beslutas 8
8542 beslutat 17
8543 beslutats 6
8544 besluten 29
8545 beslutet 38
8546 beslutets 1
8547 beslutna 3
8548 besluts- 2
8549 beslutsam 4
8550 beslutsamhet 17
8551 beslutsamma 1
8552 beslutsamt 10
8553 beslutscentrum 2
8554 beslutscentrumen 1
8555 beslutsfattande 22
8556 beslutsfattandet 10
8557 beslutsfattandets 1
8558 beslutsfattare 5
8559 beslutsfattarna 5
8560 beslutsfrihet 1
8561 beslutsförfaranden 1
8562 beslutsförfarandena 1
8563 beslutsförfarandet 1
8564 beslutsmakt 1
8565 beslutsmakten 2
8566 beslutsnivå 1
8567 beslutsorgan 1
8568 beslutsposter 1
8569 beslutsprocess 4
8570 beslutsprocessen 25
8571 beslutsprocesser 2
8572 beslutsprocesserna 4
8573 beslutsrätt 3
8574 beslutsstrukturer 1
8575 beslutstyperna 1
8576 beslutsunderlag 1
8577 beslutsunderlaget 2
8578 besläktade 1
8579 beslöt 13
8580 bespara 3
8581 besparade 1
8582 besparar 2
8583 besparingar 6
8584 besparings- 1
8585 best 4
8586 bestod 6
8587 bestraffa 1
8588 bestraffade 1
8589 bestraffar 2
8590 bestraffas 7
8591 bestraffning 1
8592 bestraffningar 1
8593 bestrida 4
8594 bestrider 1
8595 bestrids 2
8596 bestrålning 1
8597 bestyrka 1
8598 beställa 1
8599 beställde 2
8600 beställdes 1
8601 beställningar 2
8602 beställt 3
8603 beställts 1
8604 bestämd 7
8605 bestämda 14
8606 bestämdaste 2
8607 bestämde 6
8608 bestämdhet 2
8609 bestämma 22
8610 bestämmas 2
8611 bestämmelse 11
8612 bestämmelsen 3
8613 bestämmelsens 1
8614 bestämmelser 117
8615 bestämmelserna 57
8616 bestämmer 8
8617 bestäms 4
8618 bestämt 41
8619 bestämts 1
8620 beständig 2
8621 bestå 8
8622 bestående 14
8623 bestånd 8
8624 bestånden 8
8625 beståndet 3
8626 beståndsdel 11
8627 beståndsdelar 15
8628 beståndsdelarna 3
8629 beståndsdelen 1
8630 består 42
8631 bestått 1
8632 bestört 1
8633 bestörtning 3
8634 besudlade 2
8635 besvara 30
8636 besvarade 2
8637 besvarades 1
8638 besvarandet 1
8639 besvarar 4
8640 besvaras 9
8641 besvarat 1
8642 besvarats 2
8643 besvikelse 11
8644 besviken 9
8645 besviket 1
8646 besvikna 5
8647 besvär 2
8648 besvära 1
8649 besvärades 1
8650 besväret 3
8651 besvärlig 5
8652 besvärliga 5
8653 besvärligare 2
8654 besvärligt 2
8655 besynnerlig 2
8656 besynnerliga 2
8657 besynnerligheter 2
8658 besynnerligt 1
8659 besättning 3
8660 besättningen 2
8661 besök 29
8662 besöka 7
8663 besökare 3
8664 besökarna 1
8665 besöket 2
8666 besöksnäringens 1
8667 besökt 1
8668 besökte 6
8669 beta 1
8670 betade 1
8671 betala 83
8672 betalade 5
8673 betalar 48
8674 betalas 6
8675 betalat 6
8676 betalats 7
8677 betalbara 1
8678 betalbart 1
8679 betald 1
8680 betalda 2
8681 betalning 2
8682 betalningar 6
8683 betalningen 1
8684 betalningsansvariga 1
8685 betalningsbemyndiganden 1
8686 betalningsförmågan 1
8687 betalningsförseningar 1
8688 betalningsmedel 1
8689 betalningsskyldiges 1
8690 betalningssystemen 1
8691 betalt 5
8692 betalts 1
8693 bete 1
8694 beteckna 3
8695 betecknade 1
8696 betecknande 2
8697 betecknar 2
8698 betecknas 5
8699 beteckningen 3
8700 betedde 1
8701 beteende 4
8702 beteendemönster 1
8703 beteenden 1
8704 beter 1
8705 betingad 1
8706 betingade 1
8707 betingar 1
8708 betingat 1
8709 betingelser 3
8710 betingelserna 1
8711 betitlat 1
8712 betjäna 3
8713 betjänas 1
8714 betjänta 1
8715 betona 68
8716 betonade 11
8717 betonades 2
8718 betonandet 1
8719 betonar 27
8720 betonas 18
8721 betonat 10
8722 betonats 1
8723 betoning 5
8724 betoningen 1
8725 betrakta 18
8726 betraktade 6
8727 betraktande 2
8728 betraktar 26
8729 betraktas 25
8730 betraktat 3
8731 betraktats 1
8732 betryggande 5
8733 beträda 1
8734 beträffade 1
8735 beträffande 68
8736 beträffar 94
8737 bett 13
8738 betungande 3
8739 betvivla 2
8740 betvivlade 1
8741 betvivlar 9
8742 betyda 7
8743 betydande 68
8744 betydde 6
8745 betydelse 146
8746 betydelsefull 11
8747 betydelsefulla 16
8748 betydelsefullt 17
8749 betydelselös 1
8750 betydelselöst 2
8751 betydelsen 29
8752 betyder 61
8753 betydligt 33
8754 betyg 1
8755 betygar 1
8756 betänk 1
8757 betänka 5
8758 betänkande 382
8759 betänkanden 25
8760 betänkandena 5
8761 betänkandet 198
8762 betänkandets 4
8763 betänker 3
8764 betänkligheter 8
8765 beundran 2
8766 beundrar 4
8767 beundrat 2
8768 bevaka 5
8769 bevakad 1
8770 bevakade 1
8771 bevakar 3
8772 bevakaren 1
8773 bevakning 2
8774 bevara 55
8775 bevarad 2
8776 bevarade 1
8777 bevarande 26
8778 bevarandeområde 2
8779 bevarandet 12
8780 bevarar 5
8781 bevaras 6
8782 bevarats 2
8783 bevattning 3
8784 beveka 1
8785 bevekande 1
8786 bevilja 24
8787 beviljad 1
8788 beviljade 6
8789 beviljades 1
8790 beviljande 4
8791 beviljanden 2
8792 beviljandet 4
8793 beviljar 9
8794 beviljas 12
8795 beviljat 7
8796 beviljats 8
8797 bevis 53
8798 bevisa 14
8799 bevisad 1
8800 bevisade 1
8801 bevisades 1
8802 bevisar 3
8803 bevisas 1
8804 bevisat 2
8805 bevisats 3
8806 bevisbörda 3
8807 bevisbördan 5
8808 bevisen 4
8809 beviset 3
8810 bevisningsfel 1
8811 bevista 1
8812 bevistade 1
8813 bevittna 2
8814 bevittnar 3
8815 bevittnat 2
8816 bevänt 1
8817 beväpnade 1
8818 beväpning 1
8819 bibehålla 19
8820 bibehållande 1
8821 bibehållandet 1
8822 bibehållas 3
8823 bibehållen 2
8824 bibehåller 5
8825 bibehållits 1
8826 bibehålls 4
8827 bibliotekarie 1
8828 bibliotekarien 1
8829 biblioteken 1
8830 bibliotekens 1
8831 bidade 1
8832 bidra 103
8833 bidrag 102
8834 bidragande 2
8835 bidragen 7
8836 bidraget 7
8837 bidragit 20
8838 bidragsberoende 1
8839 bidragsgivare 3
8840 bidragsgivaren 3
8841 bidragsgivarna 4
8842 bidragsgivning 1
8843 bidragshjälp 1
8844 bidragsnarkomaner 1
8845 bidrar 52
8846 bidrog 6
8847 bieffekt 1
8848 bieffekter 2
8849 bieffekterna 1
8850 bifall 7
8851 bifalla 1
8852 bifallas 3
8853 bifallit 1
8854 biff 1
8855 bifloder 1
8856 bifogade 1
8857 bifogat 1
8858 bifångster 1
8859 bifångsterna 1
8860 biföll 4
8861 big 1
8862 bigotteri 1
8863 bil 19
8864 bil- 1
8865 bilaga 6
8866 bilagan 3
8867 bilagor 1
8868 bilagorna 4
8869 bilagts 1
8870 bilar 63
8871 bilarbetare 1
8872 bilarna 8
8873 bilarnas 2
8874 bilatera 1
8875 bilateral 3
8876 bilaterala 12
8877 bilateralt 6
8878 bilbeståndet 1
8879 bilbranschen 1
8880 bild 37
8881 bilda 14
8882 bildade 3
8883 bildades 5
8884 bildande 2
8885 bildandet 8
8886 bildar 10
8887 bildas 12
8888 bildat 2
8889 bildats 2
8890 bildelar 2
8891 bildelarna 1
8892 bilden 10
8893 bilder 4
8894 bilderna 1
8895 bildligt 1
8896 bildningar 1
8897 bildnings- 1
8898 bildtext 1
8899 bildvisningsinformation 1
8900 bilen 23
8901 bilens 1
8902 bilindustri 6
8903 bilindustrin 18
8904 bilindustrins 5
8905 bilindustris 2
8906 bilister 1
8907 bilisterna 1
8908 biljetten 1
8909 biljoner 1
8910 bilkonstruktörerna 1
8911 bilkyrkogårdar 1
8912 bilköpare 2
8913 billig 1
8914 billiga 2
8915 billigare 7
8916 billigaste 1
8917 billigt 4
8918 bilmärke 1
8919 bilnyckeln 1
8920 bilolyckan 1
8921 bilpark 2
8922 bilparken 4
8923 bilpriset 1
8924 bilproduktion 1
8925 bils 2
8926 bilsektorns 1
8927 bilskrotningen 1
8928 bilskrotningsmetod 1
8929 biltillverkare 4
8930 biltillverkaren 1
8931 biltillverkares 1
8932 biltillverkarna 8
8933 biltillverkarnas 1
8934 biltillverkning 1
8935 bilvrak 4
8936 bilvraket 2
8937 bilägarna 1
8938 bilägga 1
8939 bilåtervinningsmarknaden 1
8940 bin 2
8941 binda 4
8942 bindande 35
8943 bindas 1
8944 binder 3
8945 bio 2
8946 biodiversitet 1
8947 biografi 1
8948 biologer 1
8949 biologisk 8
8950 biologiska 22
8951 biologiskt 2
8952 biomassa 1
8953 bioplast 1
8954 biosfären 1
8955 biosäkerhet 1
8956 biosäkerhetsprotokollet 1
8957 biotekniken 2
8958 biotekniska 1
8959 biotoperna 1
8960 bisarra 1
8961 bister 1
8962 bistå 7
8963 bistånd 41
8964 biståndet 10
8965 bistånds 1
8966 biståndsflödena 2
8967 biståndsfrågor 1
8968 biståndsgivare 1
8969 biståndsgivaren 4
8970 biståndshjälp 1
8971 biståndsideologin 1
8972 biståndsmottagare 1
8973 biståndspengarna 2
8974 biståndspolitik 1
8975 biståndspolitiken 1
8976 biståndsprogram 1
8977 biståndsprogrammen 2
8978 biståndssystem 1
8979 biståndsvolym 1
8980 bistår 1
8981 bistått 3
8982 bit 12
8983 bitande 1
8984 bitar 7
8985 biter 2
8986 bitmappar 1
8987 biträdande 1
8988 biträdas 1
8989 biträde 1
8990 bitter 3
8991 bitterhet 1
8992 bittert 1
8993 bitti 1
8994 bittra 1
8995 bjuda 5
8996 bjudande 1
8997 bjuder 2
8998 bjudit 2
8999 bjärt 1
9000 bjärtare 1
9001 bjöd 2
9002 björnman 1
9003 bl 3
9004 bl.a. 49
9005 blackmail 1
9006 blad 1
9007 bladen 1
9008 blamerande 1
9009 bland 162
9010 blanda 11
9011 blandad 1
9012 blandade 2
9013 blandar 5
9014 blandas 4
9015 blandat 3
9016 blandning 5
9017 blandningar 2
9018 blandningen 2
9019 blandningens 1
9020 blandskogar 1
9021 blanka 1
9022 blanketter 1
9023 blanko 1
9024 blanksteg 1
9025 blankt 1
9026 bleckhink 1
9027 bleiben 1
9028 blek 2
9029 bleka 5
9030 blekaste 1
9031 blekgult 1
9032 bleknar 1
9033 bleknat 1
9034 blekningsmedel 1
9035 blekt 1
9036 blev 111
9037 bli 424
9038 blick 17
9039 blicka 1
9040 blickar 4
9041 blickarna 1
9042 blicken 8
9043 blickfältet 1
9044 blickpunkten 1
9045 blind 5
9046 blinda 2
9047 blinka 1
9048 blinkade 6
9049 blinkar 1
9050 blint 4
9051 blir 305
9052 blivande 1
9053 blivit 107
9054 blixt 2
9055 blixtar 1
9056 blixtlås 1
9057 blixtrande 1
9058 blixtvisit 1
9059 blixtärr 1
9060 block 3
9061 blockad 3
9062 blockaden 7
9063 blockadinstrument 1
9064 blockbildning 1
9065 blockera 5
9066 blockerad 2
9067 blockerade 2
9068 blockerar 4
9069 blockeras 3
9070 blockerat 3
9071 blockering 1
9072 blocket 1
9073 blod 7
9074 blodbad 1
9075 blodet 1
9076 blodfläckad 1
9077 blodigt 2
9078 blodspillan 1
9079 blomma 2
9080 blommade 1
9081 blommig 1
9082 blommiga 1
9083 blommigt 1
9084 blommor 6
9085 blomrabatterna 1
9086 blomsternoter 1
9087 blomstrande 1
9088 blomstrar 1
9089 blomstring 2
9090 blond 3
9091 blonda 1
9092 blonde 1
9093 blont 1
9094 blott 2
9095 blotta 1
9096 blottade 1
9097 blottades 1
9098 blottas 1
9099 blunda 4
9100 blundar 4
9101 bly 5
9102 blyga 1
9103 blyghet 1
9104 blygrått 1
9105 blygsam 4
9106 blygsamhet 3
9107 blygsamma 6
9108 blygsammare 1
9109 blygsamt 2
9110 blyregnet 1
9111 bläckfläckar 1
9112 bläckställ 1
9113 bländade 1
9114 bländande 5
9115 blänka 1
9116 blänkande 1
9117 blänkte 2
9118 blå 15
9119 blåa 1
9120 blåfenad 8
9121 blåfenade 3
9122 blågrön 1
9123 blåkläder 1
9124 blåsa 1
9125 blåser 1
9126 blåslagen 1
9127 blåste 4
9128 blåstes 1
9129 blått 5
9130 blöt 2
9131 blöta 1
9132 bo 8
9133 bodde 11
9134 boende 3
9135 bogsera 2
9136 bogserade 1
9137 bogserarna 1
9138 bogserbåt 3
9139 bogserbåtar 1
9140 bojkott 1
9141 bojkotta 1
9142 bojkottar 1
9143 bojkotten 1
9144 bok 20
9145 bokad 1
9146 boken 9
9147 bokens 1
9148 bokföring 1
9149 bokföringsbegrepp 1
9150 bokhandeln 2
9151 boklista 1
9152 bokmärket 1
9153 bokslut 3
9154 bokstaven 1
9155 bokstavligen 5
9156 bokstavligt 1
9157 bokstäver 1
9158 bokstäverna 1
9159 bokälskare 1
9160 bolag 7
9161 bolagen 2
9162 bolagens 2
9163 bolaget 4
9164 bolagets 1
9165 bolags 2
9166 bolagsskatter 2
9167 bollen 3
9168 bollspel 1
9169 bolsjevikiska 1
9170 bolsjevitisk 1
9171 bomb 7
9172 bomba 1
9173 bombades 1
9174 bombardera 1
9175 bombarderade 1
9176 bombattentat 1
9177 bomben 1
9178 bomber 2
9179 bombexplosioner 1
9180 bombning 1
9181 bombningar 6
9182 bombningarna 5
9183 bombningen 1
9184 bomull 1
9185 bomullskjorta 1
9186 bomullstyger 2
9187 bon 1
9188 bondedans 1
9189 bondens 1
9190 bondgård 1
9191 bondgården 1
9192 bondkvinna 1
9193 bonus 1
9194 boom 1
9195 booming 1
9196 bor 46
9197 bord 10
9198 borde 243
9199 bordeauxvin 1
9200 borden 1
9201 bordet 9
9202 bordlades 1
9203 bords 1
9204 bordsgaffeln 1
9205 bordsgrannens 1
9206 bordstal 1
9207 borga 1
9208 borgar 2
9209 borgen 1
9210 borgenärernas 1
9211 borgerlig 1
9212 borgmästare 8
9213 borgmästarens 1
9214 borgmästarinna 1
9215 borgmästarna 1
9216 borrar 3
9217 borsta 2
9218 borstade 2
9219 borstat 1
9220 bort 137
9221 borta 13
9222 bortemot 1
9223 bortfaller 8
9224 bortfallet 2
9225 bortförd 1
9226 bortglömd 2
9227 bortglömda 3
9228 bortkastad 1
9229 bortkastat 2
9230 bortom 16
9231 bortprioriteras 1
9232 bortse 11
9233 bortser 6
9234 bortsett 8
9235 bortskämda 2
9236 bortsläppt 1
9237 bortsållningen 1
9238 borttagandet 1
9239 borttappat 1
9240 bortåt 1
9241 bosatt 1
9242 bosatta 6
9243 boskapsdöden 1
9244 boskapsinitiativ 1
9245 boskapsskötarnas 1
9246 boskapsskötsel 2
9247 boskapsuppfödarna 1
9248 bosnier 2
9249 bostad 2
9250 bostaden 1
9251 bostadshyror 1
9252 bostadsprojekt 1
9253 bostäder 7
9254 bosätta 3
9255 bosättare 1
9256 bosättningar 5
9257 bosättningarna 7
9258 bosättningsdirektiven 1
9259 bosättningsområdena 1
9260 bosättningsvillkoren 1
9261 bot 3
9262 bota 1
9263 botade 1
9264 botar 2
9265 botemedlet 2
9266 bott 2
9267 botten 21
9268 bottenlös 1
9269 bottenlösa 1
9270 bottnar 3
9271 bottnen 1
9272 bottom-up-koncept 1
9273 bovar 1
9274 boven 2
9275 boy 1
9276 bra 278
9277 bragdes 1
9278 brakade 1
9279 brand 2
9280 branden 1
9281 brandgula 1
9282 brandmän 1
9283 brandplatsen 1
9284 brann 2
9285 bransch 5
9286 branschen 6
9287 branscher 3
9288 branscherna 3
9289 brant 1
9290 branten 2
9291 brasan 3
9292 brast 5
9293 brave 1
9294 bred 22
9295 breda 17
9296 bredare 23
9297 bredast 2
9298 bredband 1
9299 bredbandsnät 1
9300 bredd 1
9301 bredda 5
9302 breddar 1
9303 bredde 2
9304 bredden 5
9305 breddgraden 1
9306 breder 1
9307 bredvid 20
9308 bretagniska 1
9309 bretonne 1
9310 bretonska 3
9311 brett 20
9312 brev 33
9313 brevbärare 1
9314 brevbäraren 7
9315 brevbärarens 1
9316 breven 1
9317 brevet 4
9318 brevinsamling 1
9319 brevlåda 1
9320 brevlådeföretag 1
9321 brevutbärning 1
9322 brevväxlingen 1
9323 bricka 2
9324 brickan 2
9325 brickorna 2
9326 briefing-PM 1
9327 brigad 1
9328 briljera 1
9329 brillorna 1
9330 bringa 6
9331 bringan 1
9332 bringar 1
9333 bringas 1
9334 bringat 1
9335 brinna 1
9336 brinnande 1
9337 brinner 1
9338 bris 1
9339 briserande 1
9340 briserat 1
9341 brist 56
9342 brista 1
9343 bristande 24
9344 bristen 42
9345 brister 42
9346 bristerna 10
9347 bristfällig 5
9348 bristfälliga 6
9349 bristfälligt 4
9350 brits 1
9351 britter 2
9352 brittisk 5
9353 brittiska 37
9354 brittiske 1
9355 brittiskt 4
9356 bro 5
9357 broar 4
9358 broder 1
9359 broderade 1
9360 broders 1
9361 broderskap 4
9362 broförbindelse 1
9363 brohuvuden 1
9364 brokig 1
9365 brokigt 1
9366 bromerade 5
9367 broms 1
9368 bromsa 5
9369 bromsar 4
9370 bromsas 1
9371 bromsat 1
9372 bromsen 1
9373 bromsvätska 1
9374 bronsmynten 1
9375 bror 4
9376 broregioner 1
9377 brorsdotter 1
9378 brorson 1
9379 broskbemängda 1
9380 brother 1
9381 brott 56
9382 brottas 2
9383 brottats 2
9384 brotten 2
9385 brottmål 15
9386 brottmålsdomstol 1
9387 brottmålsdomstolar 1
9388 brottmålsdomstolen 3
9389 brottningsmatchen 1
9390 brottsanklagar 1
9391 brottsbekämpning 3
9392 brottsbekämpningen 2
9393 brottsfrågor 1
9394 brottsförebyggande 1
9395 brottslig 1
9396 brottsliga 4
9397 brottslighet 9
9398 brottsligheten 15
9399 brottsling 1
9400 brottslingar 5
9401 brottslingarna 2
9402 brottsmålssidan 1
9403 brottsoffer 2
9404 brottsrubriker 1
9405 brottsskolor 1
9406 brotullarna 1
9407 bruk 14
9408 brukade 29
9409 brukar 8
9410 brukarna 1
9411 brukas 1
9412 bruket 7
9413 brummade 2
9414 brun 1
9415 bruna 5
9416 brunn 1
9417 brunnen 1
9418 brunrosa 1
9419 brunt 1
9420 brusande 1
9421 bruset 1
9422 brutal 2
9423 brutala 4
9424 brutalt 2
9425 brutit 5
9426 brutits 3
9427 bruttoinvesteringar 1
9428 bruttonationalinkomsten 3
9429 bruttonationalprodukt 2
9430 bruttonationalprodukten 2
9431 bry 5
9432 brydde 4
9433 brygga 1
9434 bryggan 1
9435 brynet 1
9436 bryr 13
9437 brysk 1
9438 bryta 16
9439 brytas 2
9440 bryter 18
9441 brytning 4
9442 brytningar 1
9443 brytningen 2
9444 brytningsåret 1
9445 bryts 1
9446 brytt 1
9447 bräcklig 2
9448 bräckliga 4
9449 bräm 1
9450 brända 2
9451 brände 2
9452 bränder 1
9453 bränderna 1
9454 bränna 3
9455 brännande 1
9456 brännas 1
9457 bränning 2
9458 bränningar 1
9459 bränningarna 1
9460 bränningen 1
9461 brännmärka 1
9462 bränsle 3
9463 bränsleförvaring 1
9464 bränslekvaliteten 1
9465 bränslen 3
9466 bränsleskatt 1
9467 bränslesnåla 2
9468 bränslesnålare 2
9469 bränslet 1
9470 bränsletransporter 1
9471 bränts 1
9472 bräsch 1
9473 bräschen 2
9474 brådska 5
9475 brådskande 46
9476 brådskar 2
9477 bråk 1
9478 bråkade 1
9479 bråkdel 2
9480 bråkdels 1
9481 bråket 1
9482 bråkiga 1
9483 bröd 6
9484 bröder 1
9485 brödskiva 1
9486 brödsäd 1
9487 bröllopet 1
9488 bröllopsnatten 1
9489 bröst 6
9490 bröstben 1
9491 brösten 2
9492 bröstet 1
9493 brösttoner 1
9494 bröt 6
9495 bröts 1
9496 bubbla 1
9497 bubblan 2
9498 bubblor 1
9499 bucklade 1
9500 buddha 1
9501 buddhistiska 1
9502 budfirmor 1
9503 budget 52
9504 budgetanslag 4
9505 budgetanslaget 1
9506 budgetanspråk 1
9507 budgetar 6
9508 budgetarbetet 1
9509 budgetarna 1
9510 budgetbalans 1
9511 budgetbehov 1
9512 budgetbeloppet 1
9513 budgetberäkning 1
9514 budgetberäkningen 1
9515 budgetbeslut 1
9516 budgetbestämmelserna 1
9517 budgetchefen 1
9518 budgetdiskussioner 1
9519 budgeteffekten 1
9520 budgeten 53
9521 budgetenhet 1
9522 budgetens 1
9523 budgetera 1
9524 budgetfråga 1
9525 budgetfrågan 3
9526 budgetfrågor 1
9527 budgetförfarande 1
9528 budgetförfarandet 2
9529 budgetförordning 2
9530 budgetförordningen 8
9531 budgetförslag 1
9532 budgetförslaget 2
9533 budgetförvaltning 2
9534 budgetgest 1
9535 budgetkonsekvenser 2
9536 budgetkontroll 1
9537 budgetkontrollen 1
9538 budgetkontrollutskott 1
9539 budgetkontrollutskottet 14
9540 budgetkontrollutskottets 1
9541 budgetkravet 1
9542 budgetmyndigheten 2
9543 budgetmässiga 2
9544 budgetnivå 1
9545 budgetnärmanden 1
9546 budgetområde 1
9547 budgetplan 6
9548 budgetplanen 9
9549 budgetplaner 1
9550 budgetplanerna 3
9551 budgetpolitik 5
9552 budgetpolitiken 1
9553 budgetpost 13
9554 budgetposten 7
9555 budgetposter 5
9556 budgetposterna 2
9557 budgetreform 1
9558 budgetrubrik 3
9559 budgetrubriker 1
9560 budgetsituation 1
9561 budgetstöd 1
9562 budgetstödet 1
9563 budgetsynpunkt 1
9564 budgetunderskott 1
9565 budgetutskott 1
9566 budgetutskottet 10
9567 budgetåret 13
9568 budgetårets 1
9569 budgetåtgärder 1
9570 budgetöverbud 1
9571 budgetöverenskommelse 1
9572 budgetövervakare 1
9573 budord 1
9574 budordet 1
9575 buds 2
9576 budskap 23
9577 budskapet 5
9578 bugade 1
9579 building 1
9580 buk 1
9581 bukiga 1
9582 bukt 2
9583 bukter 1
9584 bullar 2
9585 bulldog 1
9586 bulldozrar 1
9587 bulle 1
9588 buller 1
9589 bullgroda 1
9590 bullrigare 1
9591 bultade 2
9592 bulten 1
9593 bunden 3
9594 bundit 1
9595 bundna 1
9596 bundsförvant 1
9597 buntar 1
9598 bur 6
9599 burden 1
9600 buren 2
9601 burens 1
9602 burit 6
9603 burken 1
9604 burklocket 1
9605 burktomater 1
9606 busflin 1
9607 bushen 4
9608 business 1
9609 business-toppmötet 1
9610 buskagen 1
9611 buskar 1
9612 busken 2
9613 buskiga 1
9614 buskvegetationen 1
9615 buss 4
9616 bussar 2
9617 bussfilerna 1
9618 busslinjer 1
9619 busstjänst 1
9620 but 1
9621 buta-trä 1
9622 butelj 1
9623 butik 2
9624 butiken 4
9625 butiker 2
9626 butiksdisk 1
9627 butiksdörren 1
9628 butiksfönster 1
9629 butiksfönstren 1
9630 butiksfönstret 1
9631 butiksförsäljningen 1
9632 buttert 1
9633 buxbomsbord 1
9634 bwana 1
9635 by 6
9636 byar 3
9637 byarna 3
9638 bygga 64
9639 byggande 3
9640 byggandet 6
9641 byggas 12
9642 byggd 3
9643 byggde 3
9644 byggdes 2
9645 bygge 2
9646 bygger 24
9647 bygget 5
9648 byggets 2
9649 bygglåda 1
9650 byggmästare 1
9651 byggnad 10
9652 byggnaden 8
9653 byggnader 1
9654 byggnaderna 1
9655 byggnadstillstånd 1
9656 byggnadstillståndet 1
9657 byggs 6
9658 byggstenarna 1
9659 byggt 10
9660 byggts 3
9661 bylte 1
9662 byn 4
9663 byrå 3
9664 byråer 6
9665 byråerna 1
9666 byråkrater 1
9667 byråkraternas 1
9668 byråkrati 23
9669 byråkratin 4
9670 byråkratisk 5
9671 byråkratiska 11
9672 byråkratiskt 4
9673 byrån 5
9674 byråns 1
9675 byta 11
9676 byte 2
9677 byten 1
9678 byter 2
9679 byteshandel 1
9680 bytet 1
9681 bytts 1
9682 byxfickorna 1
9683 byxor 2
9684 byxorna 1
9685 bädd 1
9686 bägare 2
9687 bägaren 1
9688 bägge 5
9689 bälte 1
9690 bände 1
9691 bänk 2
9692 bänkarna 1
9693 bär 38
9694 bära 20
9695 bärande 3
9696 bärare 2
9697 bäras 5
9698 bärighet 1
9699 bärkraft 1
9700 bärs 3
9701 bäst 28
9702 bästa 126
9703 bäste 5
9704 bättra 1
9705 bättre 266
9706 båda 108
9707 bådadera 1
9708 både 188
9709 bågnat 1
9710 bålen 1
9711 bålrullningar 1
9712 bården 1
9713 bås 1
9714 båt 4
9715 båtar 16
9716 båtarna 4
9717 båtarnas 1
9718 båtars 1
9719 båten 1
9720 båtens 2
9721 bébé 1
9722 böcker 15
9723 böckerna 1
9724 böckling 2
9725 böcklingar 2
9726 bödelsdräng 1
9727 böja 1
9728 böjd 2
9729 böjda 1
9730 böjde 7
9731 böjelse 1
9732 böjt 1
9733 bölande 1
9734 böljande 1
9735 bön 1
9736 bönbok 1
9737 bönder 3
9738 bönderna 2
9739 bönen 1
9740 bönens 1
9741 bör 614
9742 börda 4
9743 bördan 8
9744 bördor 1
9745 bördorna 3
9746 börja 126
9747 började 64
9748 början 82
9749 börjar 59
9750 börjat 36
9751 börsen 2
9752 börser 1
9753 börsindex 1
9754 börsmarknaderna 1
9755 börsnoterade 1
9756 börsvärde 2
9757 bössan 1
9758 böter 5
9759 bötesstraff 2
9760 c 2
9761 c'est 1
9762 ca 6
9763 calendas 1
9764 calvinistiska 1
9765 can 1
9766 canapéer 1
9767 canapérecept 1
9768 cancer 2
9769 cancerböld 1
9770 cancerframkallande 1
9771 cannabisen 1
9772 capita 14
9773 caracoling 1
9774 case 1
9775 casually 1
9776 caulerpa 1
9777 cell 2
9778 celler 1
9779 celsius 1
9780 cementerar 2
9781 censurera 1
9782 cent 1
9783 centimeter 4
9784 centra 3
9785 central 29
9786 central- 3
9787 centrala 37
9788 centralafrikanska 1
9789 centralatlanten 1
9790 centralbanken 11
9791 centralbankens 4
9792 centralbanker 1
9793 centralbankerna 1
9794 centraleuropeiska 2
9795 centralförvaltningars 1
9796 centralförvaltningen 1
9797 centralisera 1
9798 centraliserad 2
9799 centraliserade 1
9800 centraliserande 1
9801 centraliserar 2
9802 centraliserat 2
9803 centraliserats 1
9804 centralisering 6
9805 centralistiska 1
9806 centralistiskt 2
9807 centralregering 2
9808 centralregeringen 2
9809 centralstyrningen 1
9810 centralt 10
9811 centre 1
9812 centrerats 1
9813 centrum 28
9814 centrumen 3
9815 ceremonier 1
9816 ceremonin 3
9817 certifiering 1
9818 certifieringssällskap 1
9819 certifikat 3
9820 champagne 3
9821 champagneflaska 1
9822 change 1
9823 chans 31
9824 chansen 7
9825 chanser 6
9826 chanserna 2
9827 chapeau 1
9828 charaderna 1
9829 charm 1
9830 charmanta 1
9831 charmen 1
9832 chartrar 1
9833 chassid 2
9834 chassiden 3
9835 chassider 2
9836 chassiderna 3
9837 chassidim 1
9838 chassidisk 1
9839 chaufförer 3
9840 check 1
9841 checken 5
9842 chef 8
9843 chefen 3
9844 chefer 5
9845 cheferna 6
9846 chefs- 1
9847 chefsjobb 1
9848 chefsrevisor 1
9849 chefstjänster 1
9850 chilenska 1
9851 chock 2
9852 chockad 2
9853 chockade 1
9854 chocken 3
9855 chocker 1
9856 chockerad 1
9857 chockerade 2
9858 chockerande 4
9859 chockerar 1
9860 chockerna 1
9861 choklad 4
9862 chokladdirektivet 1
9863 chokladvaror 1
9864 cigarett 4
9865 cigaretten 1
9866 cigaretter 2
9867 cigarettföretagets 1
9868 cigarettmärke 1
9869 cigarettpapper 1
9870 cigarettröken 1
9871 cigarr 1
9872 cigarrask 1
9873 cigarrer 1
9874 cirka 25
9875 cirkel 2
9876 cirkeldiagram 1
9877 cirkelns 1
9878 cirklar 2
9879 cirkulera 1
9880 cirkulerar 5
9881 cirkulerat 1
9882 cirkulärbrev 1
9883 citat 3
9884 citera 10
9885 citerade 1
9886 citerar 21
9887 citeras 3
9888 citrusfrukter 1
9889 civil 7
9890 civil- 1
9891 civila 52
9892 civilbefolkningen 3
9893 civilförsvaret 1
9894 civilförsvarsmakt 1
9895 civilisation 4
9896 civilisationen 1
9897 civilisationens 1
9898 civilisera 1
9899 civiliserad 4
9900 civiliserade 3
9901 civiliserat 4
9902 civilist 1
9903 civilmål 1
9904 civilperson 1
9905 civilpolis 1
9906 civilrätt 1
9907 civilrättens 1
9908 civilrättsligt 1
9909 civilskydd 2
9910 civilskyddet 1
9911 civilt 4
9912 clauses 1
9913 clearingorganisationer 1
9914 close 1
9915 clowneri 1
9916 coccidiostatika 2
9917 cocktailbjudningar 1
9918 cocktailklänning 1
9919 collage 1
9920 cologne 1
9921 combattant 1
9922 comitology 2
9923 commitment 2
9924 common 1
9925 compassion 1
9926 compounder 1
9927 con 1
9928 conditio 2
9929 conduite 1
9930 conference 1
9931 confidence 1
9932 coniuntis 1
9933 consentiment 1
9934 contradictio 1
9935 contrario 1
9936 contre-filet 1
9937 control 2
9938 controlto 1
9939 cool 1
9940 copyright 1
9941 corporate 3
9942 corpus 6
9943 correcta 2
9944 correctness 1
9945 cost-benefit-analys 5
9946 costing 1
9947 counter 1
9948 counter-instrument 1
9949 countries 1
9950 coup 1
9951 cowboy 2
9952 cowboystövlar 1
9953 creams 1
9954 crescendo 1
9955 cricketmatcher 1
9956 crisis 1
9957 cyanid 3
9958 cyanidförgiftat 1
9959 cyanidtillverkning 1
9960 cyberspace 1
9961 cykel 1
9962 cykeln 1
9963 cyklade 1
9964 cyklar 1
9965 cyklonen 1
9966 cynisk 1
9967 cynism 1
9968 cypresser 1
9969 cyprioter 2
9970 cyprioterna 2
9971 cypriotiska 13
9972 cypriots 1
9973 d 2
9974 d'Enghiens 1
9975 d'argent 1
9976 d'essai 1
9977 d'etat 1
9978 d'intention 1
9979 da 9
9980 dag 592
9981 dagar 51
9982 dagarna 24
9983 dagarnas 1
9984 dagars 2
9985 dagen 27
9986 dagens 54
9987 daghemsplatser 1
9988 daglig 2
9989 dagliga 16
9990 dagligen 12
9991 dagligt 1
9992 daglönare 1
9993 dagmamma 1
9994 dagordning 43
9995 dagordningen 56
9996 dagordningens 1
9997 dagordnings 1
9998 dagosens 1
9999 dags 40
10000 dagsläget 4
10001 dagstidning 2
10002 dagstidningar 2
10003 dagstidningen 1
10004 dal 1
10005 dalen 2
10006 dalens 2
10007 dam 1
10008 damen 1
10009 damer 84
10010 damerna 1
10011 damm 10
10012 dammar 5
10013 dammen 2
10014 dammens 1
10015 dammet 1
10016 dammiga 3
10017 dams 1
10018 dans 3
10019 dansa 2
10020 dansade 2
10021 dansande 1
10022 dansar 2
10023 dansare 1
10024 dansarna 2
10025 dansat 1
10026 dansgolvet 1
10027 dansk 5
10028 danska 36
10029 danslektionerna 1
10030 dar 4
10031 darrade 3
10032 dass 1
10033 dasset 1
10034 data 68
10035 data- 1
10036 databas 4
10037 databasen 4
10038 databasens 1
10039 databaser 5
10040 databasfönstret 3
10041 databasobjekt 2
10042 datablad 8
10043 databladet 2
10044 datadelen 1
10045 dataelement 4
10046 dataexperter 1
10047 datafiler 1
10048 dataformat 3
10049 datakälla 5
10050 datakällan 3
10051 datamodellen 1
10052 datan 1
10053 dataområdet 2
10054 dataschemat 1
10055 dataskydd 1
10056 datastrukturen 3
10057 datastrukturer 1
10058 datasäkerhetsrättsligt 1
10059 datatypen 1
10060 datatyper 2
10061 datautbytesformat 1
10062 datautrustning 1
10063 datavärden 1
10064 dataåtkomstsida 16
10065 dataåtkomstsidan 4
10066 dataåtkomstsidor 3
10067 dataöverföringen 1
10068 daterad 1
10069 dato 1
10070 dator 5
10071 datorbrottslighet 1
10072 datorer 2
10073 datorisering 1
10074 datorn 5
10075 datornät 1
10076 datorskrot 1
10077 datum 21
10078 datumet 4
10079 datumvärden 1
10080 de 5840
10081 deadline 1
10082 dealt 2
10083 debatt 208
10084 debatten 190
10085 debattens 2
10086 debatter 18
10087 debattera 16
10088 debatterade 4
10089 debatterar 5
10090 debatteras 11
10091 debatterat 4
10092 debatterats 1
10093 debatterna 6
10094 debattinnehållet 2
10095 debattkväll 1
10096 debattskyldigheten 1
10097 debattunderlag 1
10098 debiteras 1
10099 debiterats 1
10100 december 46
10101 december- 1
10102 decemberveckan 1
10103 decennier 9
10104 decennierna 6
10105 decenniers 2
10106 decenniet 5
10107 decennium 7
10108 decentralisera 1
10109 decentraliserad 3
10110 decentraliserade 3
10111 decentraliserar 2
10112 decentraliseras 3
10113 decentraliserat 4
10114 decentralisering 9
10115 decentraliseringen 1
10116 decentraliseringsprocessen 1
10117 decentralistisk 1
10118 definiera 21
10119 definierad 2
10120 definierade 7
10121 definierades 2
10122 definierar 6
10123 definieras 8
10124 definierat 4
10125 definierats 2
10126 definition 24
10127 definitionen 12
10128 definitioner 5
10129 definitionerna 4
10130 definitionsmässigt 5
10131 definitiv 5
10132 definitiva 4
10133 definitivt 18
10134 deformerad 1
10135 deformitet 1
10136 degenererar 1
10137 degraderas 3
10138 deklaration 1
10139 deklarationen 1
10140 deklarera 1
10141 deklarerad 1
10142 deklarerar 1
10143 deklareras 1
10144 deklarerats 1
10145 dekor 2
10146 del 391
10147 dela 23
10148 delad 3
10149 delade 9
10150 delades 2
10151 delaktig 3
10152 delaktiga 11
10153 delaktighet 11
10154 delaktigheten 2
10155 delaktigt 2
10156 delar 134
10157 delarna 10
10158 delas 17
10159 delaspekt 1
10160 delat 8
10161 delats 15
10162 delayed 2
10163 delegater 1
10164 delegaterna 2
10165 delegation 22
10166 delegationen 19
10167 delegationens 2
10168 delegationer 4
10169 delegationerna 2
10170 delegations 1
10171 delegera 2
10172 delegeras 3
10173 delegerats 1
10174 delegering 5
10175 delegeringsartikeln 1
10176 delen 79
10177 delfiner 1
10178 delfrågor 1
10179 delgivning 1
10180 delikat 2
10181 dellösning 1
10182 delmängd 2
10183 delmål 1
10184 delning 7
10185 delprivatiseringar 1
10186 delrapporten 1
10187 dels 30
10188 delsession 1
10189 delstater 1
10190 delstaterna 1
10191 delstatsbanker 2
10192 delta 72
10193 deltaga 1
10194 deltagande 74
10195 deltagandet 2
10196 deltagare 4
10197 deltagarinriktade 1
10198 deltagarna 3
10199 deltagarnas 2
10200 deltagit 11
10201 deltar 34
10202 deltid 1
10203 deltidsarbetandets 1
10204 deltidsarbeten 1
10205 deltidssysselsättning 1
10206 deltog 12
10207 delutbetalningen 2
10208 delvis 39
10209 delägarna 1
10210 dem 641
10211 demagoger 1
10212 demagogi 6
10213 demagogiska 1
10214 demaskeras 1
10215 dementera 1
10216 dementerade 1
10217 demilitariseras 1
10218 demilitariseringen 1
10219 demografin 1
10220 demografiska 10
10221 demokrat 5
10222 demokrater 5
10223 demokraterna 1
10224 demokrati 71
10225 demokratier 1
10226 demokratierna 3
10227 demokratiernas 1
10228 demokratifråga 1
10229 demokratin 36
10230 demokratins 8
10231 demokratireform 1
10232 demokratisera 3
10233 demokratisering 3
10234 demokratiseringen 1
10235 demokratiseringens 1
10236 demokratiseringsprocesserna 1
10237 demokratisk 39
10238 demokratiska 102
10239 demokratiskt 40
10240 demonisk 1
10241 demoniskt 1
10242 demonstration 7
10243 demonstrationer 4
10244 demonstrationsprojekt 1
10245 demonstrera 3
10246 demonstrerar 1
10247 demonstrerat 1
10248 demontera 2
10249 demontering 3
10250 demonteringen 1
10251 demonteringskraven 1
10252 demonteringsverksamheten 1
10253 demoraliseringen 1
10254 den 6104
10255 denied 2
10256 denna 1358
10257 denne 16
10258 dennes 8
10259 densamma 9
10260 densamme 1
10261 departement 3
10262 departementen 5
10263 departementet 2
10264 departementsnivå 1
10265 dependent 1
10266 deponera 1
10267 deponerat 1
10268 deporteringarna 1
10269 depositioner 2
10270 der 9
10271 deras 291
10272 derivat 11
10273 derivaten 2
10274 derivatinstrument 4
10275 derivatives 1
10276 derivatprodukter 1
10277 derivatregleringen 1
10278 des 3
10279 desamma 4
10280 desertering 1
10281 desertörer 1
10282 design 2
10283 designläge 3
10284 designläget 2
10285 designmiljöer 1
10286 designsmiljö 1
10287 desinfektionsmedel 1
10288 desinfektionsmedlet 1
10289 desinficering 1
10290 desperat 8
10291 desperata 3
10292 desperation 1
10293 despoter 1
10294 despotiska 1
10295 dess 270
10296 dessa 951
10297 dessutom 99
10298 dessvärre 9
10299 destabilisera 4
10300 destabiliserande 2
10301 destilleringssamhälle 1
10302 desto 24
10303 destruktiv 2
10304 destruktiva 1
10305 det 9877
10306 detalj 12
10307 detaljanalys 1
10308 detaljbestämmelser 1
10309 detaljdata 3
10310 detaljen 1
10311 detaljer 16
10312 detaljerad 10
10313 detaljerade 16
10314 detaljerat 8
10315 detaljerna 9
10316 detaljflödet 1
10317 detaljfält 1
10318 detaljfälten 1
10319 detaljhandeln 1
10320 detaljkontroll 2
10321 detaljområden 2
10322 detaljområdet 4
10323 detaljplanet 1
10324 detaljproblem 1
10325 detaljreglerade 1
10326 detaljreglering 1
10327 detaljstyr 1
10328 detektiv 3
10329 detektivarbete 1
10330 detektivromaner 1
10331 detektivverksamhet 1
10332 detektorer 1
10333 detonation 1
10334 detsamma 26
10335 detta 2198
10336 det­ 1
10337 devalvering 1
10338 deve 1
10339 development 1
10340 di 1
10341 diagnos 1
10342 diagnosen 1
10343 diagnostik 1
10344 diagram 3
10345 diagrammet 1
10346 diagrammets 1
10347 diagramtyp 1
10348 dialog 66
10349 dialogen 35
10350 dialogens 2
10351 dialoger 1
10352 dialogerna 1
10353 dialogform 1
10354 dialogrutan 4
10355 diamant 1
10356 diamanter 1
10357 diamanterna 2
10358 die 2
10359 diektivförslaget 1
10360 diesel 2
10361 differentierad 3
10362 differentierade 1
10363 differentieras 1
10364 differentierat 1
10365 differentiering 5
10366 differentieringen 2
10367 diffusa 4
10368 différence 1
10369 dig 56
10370 digital 2
10371 digitala 7
10372 dignitären 1
10373 diken 1
10374 dikt 1
10375 diktatorer 2
10376 diktatoriska 1
10377 diktatorlärling 1
10378 diktatur 7
10379 diktaturen 2
10380 diktaturer 2
10381 diktaturerna 1
10382 dikter 2
10383 dikterade 1
10384 dikterar 1
10385 dikteras 1
10386 dikterats 1
10387 diktsamlingar 1
10388 dilemma 3
10389 dilemman 1
10390 dilettanteri 1
10391 dill 1
10392 dillkvist 1
10393 dimension 22
10394 dimensionen 16
10395 dimensioner 4
10396 dimensionerna 2
10397 dimma 6
10398 dimman 1
10399 din 13
10400 dina 8
10401 dinehbefolkningen 1
10402 dinehindianerna 4
10403 dinehindianernas 1
10404 dinglade 2
10405 dinglande 1
10406 dioxiderna 1
10407 dioxin 3
10408 dioxinkrisen 2
10409 dioxinskandalen 1
10410 dioxinskräckhistorien 1
10411 dioxinskräckupplevelsen 1
10412 diplomatbeskickningar 1
10413 diplomater 2
10414 diplomati 4
10415 diplomatin 1
10416 diplomatins 1
10417 diplomatisk 5
10418 diplomatiska 13
10419 diplomatiskt 3
10420 diplomatkår 1
10421 direct 1
10422 direkt 114
10423 direkta 17
10424 direktbeskattning 1
10425 direktdialog 2
10426 direktfinansiera 1
10427 direkthjälpen 1
10428 direktinvesteringar 1
10429 direktiv 244
10430 direktiven 16
10431 direktivens 1
10432 direktivet 173
10433 direktivets 16
10434 direktivförslag 2
10435 direktivförslaget 4
10436 direktivtext 1
10437 direktkontakt 1
10438 direktkontakten 1
10439 direktorat 3
10440 direktreaktion 1
10441 direktreklam 3
10442 direktsändes 1
10443 direktsänds 1
10444 direktör 2
10445 direktören 4
10446 direktörens 1
10447 direktörerna 1
10448 direktörstyper 1
10449 dirigera 1
10450 dirigism 1
10451 dis 1
10452 disciplin 9
10453 disciplinerade 1
10454 disciplinering 2
10455 disciplinerna 1
10456 disciplinfrågor 1
10457 disciplinråden 1
10458 disciplinära 4
10459 diset 1
10460 disk 1
10461 diska 1
10462 diskbänken 1
10463 disken 5
10464 diskho 1
10465 diskret 3
10466 diskreta 1
10467 diskretion 1
10468 diskriminera 1
10469 diskriminerade 3
10470 diskriminerande 4
10471 diskrimineras 1
10472 diskriminering 59
10473 diskrimineringar 2
10474 diskrimineringen 3
10475 diskrimineringsförslag 1
10476 diskrimineringskategori 1
10477 diskrimineringskategorierna 1
10478 diskursen 1
10479 diskussion 50
10480 diskussionen 37
10481 diskussioner 47
10482 diskussionerna 13
10483 diskussions- 1
10484 diskussionsdokument 1
10485 diskussionsforum 1
10486 diskussionsgrupp 1
10487 diskussionsprocess 1
10488 diskussionspunkt 1
10489 diskussionspunkten 1
10490 diskussionsunderlag 2
10491 diskussionsämne 2
10492 diskussionsämnen 1
10493 diskutabelt 2
10494 diskutabla 2
10495 diskutera 78
10496 diskuterade 16
10497 diskuterades 4
10498 diskuterar 67
10499 diskuteras 25
10500 diskuterat 20
10501 diskuterats 12
10502 dispenser 1
10503 disponerar 1
10504 disponeras 1
10505 disponibla 2
10506 dispositioner 1
10507 dispositionerna 2
10508 disproportion 1
10509 dispyt 1
10510 disrupters 1
10511 distans 2
10512 distansförhöret 1
10513 distanshandel 1
10514 distinktion 3
10515 distraherar 1
10516 distraheras 1
10517 distraktion 1
10518 distribuera 1
10519 distribuerar 2
10520 distribution 3
10521 distributionen 1
10522 distributionsnätens 1
10523 distributionssektorn 1
10524 distributörers 1
10525 distriktsdomare 1
10526 distriktskommissarien 2
10527 dit 39
10528 dithän 1
10529 dithörande 1
10530 ditt 7
10531 ditupp 1
10532 divaner 1
10533 diverse 14
10534 diversehandeln 1
10535 diversifiera 1
10536 diversifierade 1
10537 diversifierat 1
10538 diversifiering 1
10539 divisioner 1
10540 djungel 2
10541 djungeln 1
10542 djungelns 2
10543 djup 13
10544 djupa 12
10545 djupare 8
10546 djupaste 4
10547 djupet 12
10548 djupgående 14
10549 djuphavsfiske 1
10550 djupnade 3
10551 djupnande 1
10552 djupsinnighet 2
10553 djupt 27
10554 djur 16
10555 djur- 5
10556 djurarter 2
10557 djuren 3
10558 djurens 6
10559 djuret 2
10560 djurfoder 25
10561 djurfoderblandningar 1
10562 djurfoderbranschen 1
10563 djurfoderindustrins 1
10564 djurfoderproducenterna 1
10565 djurfodret 3
10566 djurhälsovillkor 1
10567 djurhållningen 1
10568 djurliv 2
10569 djurlivet 1
10570 djurläkemedel 1
10571 djurs 2
10572 djurskyddskriterierna 1
10573 djärv 3
10574 djärva 5
10575 djärvare 2
10576 djärvhet 2
10577 djärvt 2
10578 djävlar 1
10579 djävlarna 1
10580 djävul 4
10581 djävulen 1
10582 djävulens 1
10583 djävulska 1
10584 dock 269
10585 dockor 2
10586 dodderer 1
10587 doft 3
10588 doftande 2
10589 doftar 1
10590 doften 2
10591 dog 15
10592 dogm 1
10593 dogmatiska 1
10594 dogmen 1
10595 doktor 1
10596 doktrin 4
10597 doktrinen 1
10598 dokument 102
10599 dokumentation 1
10600 dokumentationen 1
10601 dokumenten 8
10602 dokumenterade 1
10603 dokumentet 18
10604 dokumentets 1
10605 dokumentkategorier 1
10606 dokumentskåp 1
10607 dold 3
10608 dolda 3
10609 dollar 20
10610 dollarn 3
10611 dollartecken 1
10612 dolomiten 1
10613 dolt 3
10614 dolts 1
10615 dom 20
10616 domar 9
10617 domare 11
10618 domaren 2
10619 domarkollegier 1
10620 domarna 7
10621 domarnas 1
10622 domen 3
10623 dominans 3
10624 dominansen 1
10625 dominera 3
10626 dominerades 1
10627 dominerande 12
10628 dominerar 1
10629 domineras 4
10630 domino 1
10631 dominospel 1
10632 domkretsar 1
10633 domslut 3
10634 domsrätt 1
10635 domsrätten 1
10636 domstol 13
10637 domstolar 14
10638 domstolarna 11
10639 domstolars 2
10640 domstolen 24
10641 domstolens 7
10642 domstolsavgörande 1
10643 domstolsfall 1
10644 domstolsförhandlingar 2
10645 domstolsförhandlingarna 1
10646 domstolskandidat 1
10647 domstolsmyndighet 1
10648 domstolsprocessen 1
10649 domstolssystemet 2
10650 domstolstvister 1
10651 domstolsutslag 1
10652 domstolsväsen 1
10653 domäner 1
10654 donator 1
10655 donne 1
10656 donor 1
10657 dopet 1
10658 doppade 1
10659 dos 1
10660 dosis 1
10661 dossier 1
10662 dossieren 1
10663 dot.com-företag 1
10664 dotter 7
10665 dotterdirektiv 1
10666 dov 1
10667 dra 80
10668 drabba 3
10669 drabbade 44
10670 drabbades 9
10671 drabbar 13
10672 drabbas 20
10673 drabbat 11
10674 drabbats 21
10675 drack 8
10676 drag 10
10677 dragande 2
10678 dragbilen 1
10679 dragen 6
10680 draget 3
10681 draggade 1
10682 dragit 10
10683 dragits 4
10684 dragna 1
10685 dragningskraft 1
10686 dragspel 1
10687 drake 1
10688 drakgödsel 1
10689 drakonisk 1
10690 dramat 2
10691 dramatiken 1
10692 dramatiserar 1
10693 dramatisk 6
10694 dramatiska 13
10695 dramatiskt 8
10696 draperi 1
10697 draperiet 1
10698 drar 34
10699 dras 7
10700 drastisk 2
10701 drastiska 4
10702 drastiskt 8
10703 dravel 1
10704 dreglade 1
10705 dress-shirt 1
10706 drev 7
10707 drevs 3
10708 dricka 9
10709 drickande 1
10710 drickas 1
10711 drickat 1
10712 dricker 4
10713 dricks 1
10714 dricks- 1
10715 dricksvatten 10
10716 dricksvattenförsörjning 1
10717 dricksvattenförsörjningen 2
10718 dricksvattenkvalitet 1
10719 dricksvattnet 2
10720 drift 4
10721 driften 1
10722 driftiga 1
10723 driftighet 1
10724 driftsförhållanden 1
10725 driftsverksamhet 1
10726 driftsvillkoren 1
10727 driftsäkerhet 1
10728 drink 4
10729 drinken 1
10730 driva 31
10731 drivande 3
10732 drivas 3
10733 driver 16
10734 drivfjäder 1
10735 drivfjädern 1
10736 drivgarn 3
10737 driving 1
10738 drivit 2
10739 drivkraft 6
10740 drivkraften 1
10741 drivkrafter 2
10742 drivkrafterna 1
10743 drivmotor 1
10744 drivs 6
10745 drog 27
10746 drogberoende 4
10747 drogeffekter 1
10748 droger 1
10749 drogkulturen 1
10750 drogs 5
10751 droit 2
10752 droppade 1
10753 droppe 3
10754 droppen 2
10755 drottning 2
10756 drottningens 1
10757 drottninglik 1
10758 druckit 3
10759 drucknes 1
10760 drunkna 2
10761 drunknade 2
10762 drunknar 1
10763 drunknat 2
10764 dryck 1
10765 drycker 5
10766 dryckerna 1
10767 dryfta 2
10768 dryftar 2
10769 drygt 8
10770 drägligare 1
10771 drägligt 1
10772 dräkter 2
10773 drämde 1
10774 dränka 1
10775 dränkte 2
10776 dråpslag 1
10777 dröja 5
10778 dröjde 3
10779 dröjer 5
10780 dröjsmål 6
10781 dröjt 2
10782 dröm 3
10783 drömde 2
10784 drömma 3
10785 drömmande 1
10786 drömmar 3
10787 drömmen 4
10788 drömtillfälle 1
10789 du 306
10790 dualiseras 1
10791 dubbel 5
10792 dubbelbeskattning 1
10793 dubbeldörrarna 1
10794 dubbelfinansiering 1
10795 dubbelhaka 1
10796 dubbelkontrollera 1
10797 dubbelmoral 1
10798 dubbelrunda 1
10799 dubbelskrovet 2
10800 dubbelt 5
10801 dubbelväggigt 1
10802 dubbla 21
10803 dubblera 3
10804 dubblerade 1
10805 dubbleringar 1
10806 dubbleringen 1
10807 ducka 1
10808 duga 1
10809 duger 1
10810 duggades 1
10811 dugligheten 1
10812 duk 1
10813 dukade 2
10814 dukar 1
10815 dukat 1
10816 duktig 1
10817 duktiga 2
10818 duktigt 1
10819 dum 4
10820 dumhet 3
10821 dumheter 2
10822 dumpades 1
10823 dumpandet 1
10824 dumpning 9
10825 dumt 5
10826 dunans 1
10827 dunder 1
10828 dungen 1
10829 dungens 1
10830 dunkande 2
10831 dunkel 1
10832 dunkelt 1
10833 dunklet 1
10834 dunmjuka 1
10835 duns 2
10836 dures 1
10837 duschade 1
10838 dussin 3
10839 dvala 1
10840 dvs 3
10841 dvs. 126
10842 dy 1
10843 dygder 1
10844 dygn 1
10845 dygnet 2
10846 dyka 5
10847 dyker 9
10848 dykningen 1
10849 dykt 6
10850 dylika 5
10851 dylikt 1
10852 dynamik 7
10853 dynamiken 1
10854 dynamisk 9
10855 dynamiska 10
10856 dynamiskt 2
10857 dynamitladdning 1
10858 dyngbaggar 1
10859 dynggrepen 1
10860 dynghög 1
10861 dyningen 1
10862 dyr 5
10863 dyra 3
10864 dyrare 4
10865 dyraste 2
10866 dyrbar 2
10867 dyrbart 1
10868 dyrka 1
10869 dyrkan 1
10870 dyrt 5
10871 dyster 4
10872 dystert 2
10873 dystra 4
10874 däck 4
10875 däckfabrikant 1
10876 däggdjur 2
10877 dämpa 4
10878 dämpad 1
10879 dämpades 1
10880 dämpar 1
10881 dämpas 1
10882 där 940
10883 därav 7
10884 därefter 28
10885 däremellan 1
10886 däremot 39
10887 därför 514
10888 därhemma 1
10889 därhän 3
10890 däri 1
10891 däribland 15
10892 därifrån 8
10893 därigenom 33
10894 därinne 1
10895 därmed 110
10896 därnere 1
10897 däromkring 1
10898 därpå 6
10899 därtill 3
10900 därutanför 1
10901 därute 3
10902 därvid 5
10903 då 500
10904 dåd 1
10905 dådet 1
10906 dålig 15
10907 dåliga 21
10908 dåligt 21
10909 dån 1
10910 dånade 1
10911 dånande 1
10912 dånet 1
10913 dåraktiga 3
10914 dåre 2
10915 dåvarande 3
10916 défense 2
10917 démocratique 1
10918 dö 9
10919 död 27
10920 död-och-liv 1
10921 döda 28
10922 dödade 10
10923 dödades 2
10924 dödande 1
10925 dödar 6
10926 dödas 6
10927 dödat 2
10928 dödats 3
10929 döde 1
10930 döden 3
10931 dödens 3
10932 dödfödd 1
10933 dödhet 1
10934 dödliga 2
10935 dödlighet 1
10936 dödligt 1
10937 dödläge 1
10938 dödsdomen 1
10939 dödsdömd 1
10940 dödsfall 2
10941 dödsfallen 2
10942 dödsfrekvensen 1
10943 dödskallar 1
10944 dödskampen 1
10945 dödsliknande 1
10946 dödsmärkt 1
10947 dödsoffer 1
10948 dödsrikets 1
10949 dödsstraff 4
10950 dödsstraffet 8
10951 döende 2
10952 dög 1
10953 dök 15
10954 dölja 21
10955 döljer 11
10956 döljs 7
10957 döma 20
10958 dömande 1
10959 dömas 2
10960 dömd 1
10961 dömda 2
10962 dömde 2
10963 dömer 2
10964 döms 1
10965 dömts 2
10966 döpa 1
10967 döper 3
10968 döpte 1
10969 dör 13
10970 dörr 13
10971 dörrar 6
10972 dörrarna 3
10973 dörrarnas 1
10974 dörren 32
10975 dörrhandtag 1
10976 dörrklockan 1
10977 dörrvredet 1
10978 dörröppningen 2
10979 dörröverstycken 1
10980 dött 12
10981 döttrar 1
10982 döttrarna 1
10983 döva 3
10984 döve 1
10985 e 4
10986 e-Europa 3
10987 e-Europe 2
10988 e-företagande 1
10989 e-företagandet 1
10990 e-handel 1
10991 e-handeln 6
10992 e-handelsmöjligheter 1
10993 e-mail 1
10994 e-post 4
10995 e-posthastighet 1
10996 e-sidan 1
10997 e.d. 1
10998 eau 1
10999 ebben 4
11000 ebbremsa 1
11001 ecu 7
11002 ed 1
11003 eden 1
11004 effekt 29
11005 effekten 15
11006 effekter 43
11007 effekterna 30
11008 effektfull 1
11009 effektiv 77
11010 effektiva 43
11011 effektivare 34
11012 effektivaste 3
11013 effektivisera 7
11014 effektivisering 2
11015 effektivitet 33
11016 effektiviteten 17
11017 effektivitetsargument 1
11018 effektivitetskriterier 1
11019 effektivitetssprång 1
11020 effektivt 81
11021 effektstudie 1
11022 effektuera 1
11023 efter 509
11024 efter-thirst 1
11025 efterbilda 1
11026 efterbildar 1
11027 efterblivna 1
11028 efterforskningar 4
11029 efterfrågan 18
11030 efterfrågans 1
11031 efterfrågar 2
11032 efterfrågat 1
11033 efterfrågats 2
11034 efterfråge-elasticitet 2
11035 efterfrågningar 1
11036 efterföljande 4
11037 efterföljare 1
11038 efterföljarna 1
11039 eftergift 1
11040 eftergifter 5
11041 eftergivenhet 5
11042 eftergivenheten 1
11043 eftergivna 1
11044 eftergymnasial 1
11045 efterhand 11
11046 efterhandsgranskning 1
11047 efterhandskontrollen 1
11048 efterkommande 1
11049 efterkälken 3
11050 efterlevas 2
11051 efterlevnad 6
11052 efterlevs 8
11053 efterlevts 2
11054 efterlikna 2
11055 efterlysa 1
11056 efterlyser 3
11057 efterlyses 1
11058 efterlysning 1
11059 efterlyst 1
11060 efterlämnade 1
11061 eftermiddag 20
11062 eftermiddagarna 1
11063 eftermiddagen 5
11064 eftermiddagens 1
11065 eftermiddags 3
11066 eftermiddagskaffe 1
11067 eftermiddagsmyntor 1
11068 eftermiddan 1
11069 eftermäle 1
11070 efterrättstårta 1
11071 eftersatta 11
11072 eftersatthet 3
11073 eftersatthetskriteriet 1
11074 eftersläpning 4
11075 eftersläpningen 1
11076 eftersom 567
11077 eftersträva 6
11078 eftersträvade 6
11079 eftersträvansvärda 1
11080 eftersträvansvärt 1
11081 eftersträvar 9
11082 eftersträvas 5
11083 eftersträvat 1
11084 eftertanke 7
11085 eftertraktade 1
11086 eftertraktar 1
11087 eftertryck 5
11088 eftertryckligen 5
11089 efterträdare 1
11090 efterträdaren 1
11091 efterträdde 1
11092 eftertänksamhet 1
11093 efterverkningar 1
11094 efteråt 7
11095 egen 115
11096 egenansvar 1
11097 egenart 1
11098 egendom 7
11099 egendomen 1
11100 egendomlig 2
11101 egendomligheter 1
11102 egendomligt 6
11103 egendoms 1
11104 egendomsrätt 1
11105 egenföretagande 1
11106 egenföretagare 3
11107 egenföretagarna 1
11108 egenhet 2
11109 egenintresse 1
11110 egenskap 52
11111 egenskapen 11
11112 egenskaper 9
11113 egenskaperna 3
11114 egenskapsbladet 2
11115 egenskapsinställning 1
11116 egenskapsinställningar 1
11117 egenskapsinställningarna 1
11118 egenskapsinställningen 1
11119 egenskapsrutan 1
11120 egentlig 2
11121 egentliga 5
11122 egentligen 122
11123 egentligt 1
11124 egenutvecklade 1
11125 eget 77
11126 egg 1
11127 eggande 1
11128 egna 126
11129 egoism 1
11130 egoistiska 4
11131 egyptiska 3
11132 egyptiskt 1
11133 ej 40
11134 ekade 1
11135 ekologisk 8
11136 ekologiska 28
11137 ekologiskt 10
11138 ekon 1
11139 ekonom 1
11140 ekonomer 1
11141 ekonomernas 1
11142 ekonometriska 1
11143 ekonomi 92
11144 ekonomi- 2
11145 ekonomier 17
11146 ekonomierna 7
11147 ekonomiernas 1
11148 ekonomin 74
11149 ekonomins 9
11150 ekonomisk 151
11151 ekonomiska 398
11152 ekonomiske 1
11153 ekonomiskt 83
11154 ekonomiskt-finansiellt 1
11155 ekonomistyrning 9
11156 ekonomistyrningen 4
11157 ekonomisystemet 1
11158 ekosocial 1
11159 ekosystem 8
11160 ekosystemen 6
11161 ekosystemet 5
11162 ekoturism 1
11163 ekvation 1
11164 ekvatorn 1
11165 ekvilibristik 1
11166 el 1
11167 el- 3
11168 el-Sheikh 3
11169 el-Sheikh-avtalet 1
11170 elak 1
11171 elasticitet 1
11172 eld 3
11173 eldade 1
11174 elden 7
11175 eldkvast 1
11176 eldsken 1
11177 eldskenet 2
11178 eldslåga 1
11179 eldstaden 1
11180 eldsvådan 1
11181 electronic 1
11182 elefant 1
11183 elegans 1
11184 elegant 1
11185 eleganta 1
11186 elektricitet 3
11187 elektriskt 6
11188 elektrochock 1
11189 elektronik- 1
11190 elektronikavfall 1
11191 elektronikbranschen 1
11192 elektronikindustrin 1
11193 elektronisk 8
11194 elektroniska 13
11195 elektroniskt 9
11196 element 25
11197 elementet 3
11198 elementnamn 2
11199 elementära 5
11200 elevhemmets 1
11201 elfenben 4
11202 elfenbenslandet 1
11203 elfte 2
11204 eliminera 11
11205 eliminerade 1
11206 eliminerar 1
11207 elimineras 1
11208 eliminerats 1
11209 eliminering 1
11210 elit 3
11211 eliten 1
11212 elits 1
11213 elitutbildning 1
11214 elkostnaderna 1
11215 elle 1
11216 eller 1270
11217 elmaster 1
11218 eloge 2
11219 elräkningar 1
11220 elva 9
11221 elände 1
11222 eländet 1
11223 eländig 2
11224 eländiga 1
11225 emalj 1
11226 emanciperad 1
11227 embargo 2
11228 embargot 5
11229 emblem 1
11230 emblemet 1
11231 embryo 1
11232 embryoform 1
11233 embryostadiet 1
11234 emedan 1
11235 emellan 14
11236 emellanåt 3
11237 emellertid 168
11238 emigration 1
11239 emigrera 2
11240 emissionsgarantier 1
11241 emot 166
11242 emotionell 1
11243 emotionella 1
11244 emotionellt 2
11245 emotser 1
11246 empiriskt 1
11247 en 8621
11248 en-mängd 1
11249 ena 111
11250 enad 2
11251 enade 16
11252 enades 3
11253 enahanda 1
11254 enande 1
11255 enandet 2
11256 enar 1
11257 enas 9
11258 enastående 9
11259 enat 2
11260 enats 8
11261 enbart 95
11262 encefalopati 1
11263 end 1
11264 enda 191
11265 endast 217
11266 endaste 1
11267 ende 3
11268 endemisk 2
11269 endemiska 1
11270 endocrine 1
11271 endogen 1
11272 endogena 1
11273 ene 2
11274 energi 35
11275 energi- 1
11276 energiagenturer 1
11277 energianvändning 6
11278 energibesparing 3
11279 energibesparingar 1
11280 energicentra 1
11281 energidistribution 1
11282 energieffektiva 1
11283 energieffektivitet 2
11284 energier 2
11285 energierna 1
11286 energiformer 1
11287 energiförbrukningen 1
11288 energiförråden 1
11289 energiförsörjning 1
11290 energiförsörjningen 1
11291 energiförsörjningssystem 1
11292 energiimport 2
11293 energikapacitet 1
11294 energikontrollsystem 1
11295 energikrävande 1
11296 energikälla 2
11297 energikällor 34
11298 energikällorna 4
11299 energikällornas 1
11300 energimarknaden 1
11301 energimixen 1
11302 energin 4
11303 energinäten 2
11304 energiområdet 1
11305 energipolitiken 2
11306 energipotential 1
11307 energiproduktion 2
11308 energiproduktionen 1
11309 energiprogram 1
11310 energiprogrammets 1
11311 energiresurser 1
11312 energisektor 1
11313 energisektorerna 1
11314 energisektorn 4
11315 energisk 1
11316 energiska 1
11317 energiskt 4
11318 energisnåla 1
11319 energiutvinning 1
11320 energiåtervinning 1
11321 energiöverföring 1
11322 enerverande 1
11323 enes 1
11324 enfaldiga 1
11325 enformig 1
11326 enformighet 1
11327 enfranchisement 1
11328 engagemang 43
11329 engagemanget 4
11330 engagera 14
11331 engagerad 2
11332 engagerade 11
11333 engagerar 9
11334 engageras 3
11335 engagerat 4
11336 engelsk 2
11337 engelsk-franska 1
11338 engelska 29
11339 engelskspråkiga 2
11340 engelskt 2
11341 engelsman 4
11342 engelsmannen 1
11343 engelsmän 2
11344 engelsmännen 3
11345 engångsåtgärder 1
11346 enhet 19
11347 enheten 4
11348 enheter 12
11349 enheterna 6
11350 enhetlig 27
11351 enhetliga 15
11352 enhetlighet 8
11353 enhetligt 17
11354 enhetsakten 1
11355 enhetschefer 3
11356 enhetscheferna 1
11357 enhetsorganisationen 2
11358 enhetspolitiska 1
11359 enhetspris 1
11360 enhetsstat 1
11361 enhällig 3
11362 enhälliga 4
11363 enhällighet 21
11364 enhälligheten 2
11365 enhällighetsprincip 1
11366 enhällighetsprincipen 2
11367 enhälligt 28
11368 enig 2
11369 eniga 6
11370 enighet 18
11371 enigheten 1
11372 enigt 1
11373 enkel 20
11374 enkelhet 1
11375 enkelhetens 1
11376 enkelmajoritet 1
11377 enkelriktat 1
11378 enkelt 90
11379 enkelväggigt 2
11380 enkla 21
11381 enklare 8
11382 enklast 1
11383 enklaste 2
11384 enlighet 114
11385 enligt 281
11386 enmansföretag 1
11387 enorm 21
11388 enorma 50
11389 enormt 25
11390 enpartisystemet 1
11391 ens 73
11392 ensam 11
11393 ensamma 15
11394 ensamrätt 2
11395 ensamrätten 2
11396 ensamstående 2
11397 ensamt 4
11398 ense 8
11399 ensidig 4
11400 ensidiga 3
11401 ensidigt 8
11402 enskild 15
11403 enskilda 65
11404 enskildas 2
11405 enskilde 5
11406 enskildhet 1
11407 enskildheter 1
11408 enskilt 13
11409 enstaka 11
11410 entiteten 1
11411 entiteter 1
11412 entreprenad 2
11413 entreprenadföretag 1
11414 entreprenör 1
11415 entreprenören 1
11416 entreprenörerna 2
11417 entreprenörsandan 1
11418 entreprenörskap 3
11419 entreprises 2
11420 enträgen 1
11421 enträget 1
11422 entréhallen 1
11423 entusiasm 11
11424 entusiasmen 1
11425 entusiasmerande 2
11426 entusiastisk 1
11427 entusiastiskt 2
11428 entydig 1
11429 entydiga 3
11430 entydigt 6
11431 envar 1
11432 envetenheten 1
11433 envetet 1
11434 envis 1
11435 envisades 3
11436 envisas 2
11437 envishet 6
11438 envist 4
11439 enväldig 1
11440 enögd 1
11441 epidemier 3
11442 episoden 1
11443 epok 4
11444 epoken 2
11445 epokgörande 1
11446 er 571
11447 era 100
11448 erbjuda 31
11449 erbjudande 2
11450 erbjudanden 2
11451 erbjudandet 2
11452 erbjudas 3
11453 erbjuder 26
11454 erbjudit 1
11455 erbjudits 2
11456 erbjuds 6
11457 erbjöd 6
11458 erbjöds 1
11459 erfara 3
11460 erfaren 1
11461 erfarenhet 28
11462 erfarenheten 5
11463 erfarenheter 40
11464 erfarenheterna 10
11465 erfarenhetsutbyte 5
11466 erfarenhetsutbytet 2
11467 erfarit 2
11468 erfarna 1
11469 erfor 1
11470 erforderlig 3
11471 erforderliga 7
11472 erhalten 1
11473 erhålla 4
11474 erhållande 1
11475 erhåller 3
11476 erhållit 7
11477 erhållits 1
11478 erhöll 4
11479 erinra 28
11480 erinrade 7
11481 erinran 1
11482 erinrar 6
11483 erinras 2
11484 erkänd 8
11485 erkända 4
11486 erkände 6
11487 erkändes 3
11488 erkänds 1
11489 erkänna 32
11490 erkännande 31
11491 erkännandet 5
11492 erkännas 8
11493 erkänner 25
11494 erkänns 5
11495 erkänt 3
11496 erkänts 2
11497 eroderar 1
11498 ersatt 3
11499 ersatta 1
11500 ersatts 3
11501 ersätta 31
11502 ersättas 9
11503 ersätter 6
11504 ersättning 16
11505 ersättningar 4
11506 ersättningarna 1
11507 ersättningen 2
11508 ersättningsansvar 2
11509 ersättningsansvaret 1
11510 ersättningsbeloppet 1
11511 ersättningsmedel 1
11512 ersättningsnivåerna 1
11513 ersättningssystemet 1
11514 ersätts 3
11515 ert 136
11516 erövra 2
11517 erövrades 1
11518 erövrar 1
11519 erövrare 1
11520 erövring 1
11521 erövringen 1
11522 erövringståg 1
11523 es 1
11524 eskort 1
11525 eskorteras 1
11526 esogena 1
11527 esprit 1
11528 essensen 1
11529 essere 1
11530 essäer 1
11531 est 1
11532 esterno 2
11533 estetiska 1
11534 estraden 1
11535 et 3
11536 etablera 9
11537 etablerad 3
11538 etablerade 6
11539 etablerar 2
11540 etablerat 2
11541 etablerats 2
11542 etablering 3
11543 etableringskriteriet 1
11544 etablissemangets 1
11545 etapp 6
11546 etappen 4
11547 etapper 4
11548 etappvis 1
11549 etc 1
11550 etc. 11
11551 etik 1
11552 etikett 4
11553 etiketten 1
11554 etisk 1
11555 etiska 2
11556 etiskt 1
11557 etnisk 11
11558 etniska 27
11559 etniskt 8
11560 etsad 1
11561 ett 4693
11562 etthundranio 1
11563 ettåriga 1
11564 ettårsplanen 1
11565 eukalyptusträd 1
11566 euro 124
11567 euro-staterna 1
11568 euro-äventyret 1
11569 eurofederalistiska 2
11570 euron 43
11571 eurons 6
11572 euroområdet 4
11573 europaparlamentariker 2
11574 europapatent 1
11575 europatjänsteman 1
11576 europavänlig 1
11577 europeiseras 1
11578 europeisering 1
11579 europeisk 222
11580 europeiska 577
11581 europeiske 4
11582 europeiskt 62
11583 europeistisk 1
11584 europrojektet 1
11585 europé 6
11586 européen 1
11587 européer 27
11588 européerna 8
11589 européernas 3
11590 européers 2
11591 euror 2
11592 eurosedlar 1
11593 euroskeptikerna 1
11594 euroskeptiska 1
11595 eurosymboler 1
11596 eutrofiering 1
11597 evakueras 1
11598 evalueringsbefogenheter 1
11599 evenemang 2
11600 eventuell 16
11601 eventuella 32
11602 eventuellt 38
11603 evig 1
11604 eviga 3
11605 evighet 3
11606 evigt 5
11607 ex 10
11608 exakt 47
11609 exakta 17
11610 exakthet 3
11611 examen 5
11612 examensbevis 1
11613 examensbevisen 1
11614 examination 1
11615 examineringsformer 1
11616 examineringskraven 5
11617 examineringsorganen 1
11618 examineringsorganet 1
11619 examineringsvillkoren 1
11620 excellence 1
11621 exceptionell 4
11622 exceptionellt 5
11623 exempel 303
11624 exempelvis 81
11625 exemplar 8
11626 exemplarisk 1
11627 exemplariska 1
11628 exemplariskt 3
11629 exemplen 6
11630 exemplet 11
11631 exigé 1
11632 exilregeringen 1
11633 exiltibetanerna 1
11634 existens 6
11635 existensberättigande 1
11636 existensen 1
11637 existenser 2
11638 existensrätten 1
11639 existentiella 1
11640 existera 7
11641 existerade 1
11642 existerande 6
11643 existerar 27
11644 exklusiv 2
11645 exklusiva 5
11646 exklusivt 1
11647 exkrementer 1
11648 exotisk 1
11649 exotiska 1
11650 expandera 4
11651 expanderande 1
11652 expanderar 2
11653 expansion 1
11654 expansionistiska 1
11655 expansionspolitik 1
11656 expansiva 1
11657 expeditioner 1
11658 expeditionskommission 1
11659 experiment 3
11660 experimentella 1
11661 experimentera 1
11662 experimentet 1
11663 experimentroll 1
11664 experimentstadiet 2
11665 expert 1
11666 experten 1
11667 experter 15
11668 experterna 10
11669 expertgrupp 2
11670 expertgruppen 2
11671 expertgruppens 2
11672 experthjälp 1
11673 expertis 3
11674 expertkommitté 4
11675 expertkommittén 12
11676 expertkommitténs 4
11677 expertkunskap 1
11678 expertrapport 1
11679 expertregeringar 1
11680 expertutskott 1
11681 explicit 2
11682 exploatera 1
11683 exploateras 2
11684 exploaterbara 1
11685 exploatering 3
11686 exploateringen 2
11687 explodera 1
11688 exploderade 1
11689 exploderar 2
11690 explosion 3
11691 explosionen 2
11692 explosioner 1
11693 explosionsartad 1
11694 explosionsrisk 1
11695 explosiv 1
11696 exponentiell 3
11697 exponerar 1
11698 exponeras 1
11699 exponering 1
11700 export 9
11701 exportbidrag 1
11702 exportbidragen 1
11703 exportbidragssystemet 1
11704 exportbranscherna 1
11705 exporten 8
11706 exportera 14
11707 exporterar 6
11708 exporteras 4
11709 exporterat 1
11710 exporterna 1
11711 exportindustrier 1
11712 exportintäkterna 2
11713 exportkrediter 1
11714 exportkreditgarantier 1
11715 exportkreditlicens 1
11716 exportkvot 1
11717 exportör 1
11718 exportörer 2
11719 exportörerna 1
11720 expressbud 1
11721 expressfart 1
11722 expresstjänstesektorn 1
11723 extas 1
11724 extern 3
11725 externa 22
11726 externt 4
11727 extra 34
11728 extraordinär 1
11729 extraordinära 3
11730 extraordinärt 2
11731 extrarum 1
11732 extrem 1
11733 extrema 7
11734 extremhögern 10
11735 extremhögerns 6
11736 extremism 2
11737 extremistaktioner 1
11738 extremister 2
11739 extremistiska 3
11740 extremistiskt 2
11741 extremsituationer 1
11742 extremt 17
11743 f 1
11744 f.d. 20
11745 fabrik 6
11746 fabriken 6
11747 fabrikens 1
11748 fabriker 5
11749 fabrikerna 1
11750 faciliteter 1
11751 facility 1
11752 facken 1
11753 fackförbund 1
11754 fackföreningar 5
11755 fackföreningarna 4
11756 fackföreningen 1
11757 fackföreningsrörelsen 1
11758 fackföreningsrörelsens 1
11759 fackkunskaper 1
11760 facklan 1
11761 fackliga 3
11762 fackmässig 1
11763 fackrörelsen 1
11764 facktermer 1
11765 fact 1
11766 facto 2
11767 fadder 1
11768 fadern 1
11769 faders 1
11770 failures 1
11771 faire 1
11772 fakta 13
11773 faktabas 1
11774 faktainsamlingsresa 2
11775 faktaunderlag 1
11776 faktisk 3
11777 faktiska 14
11778 faktiskt 145
11779 faktor 25
11780 faktorer 30
11781 faktorerna 2
11782 faktorn 5
11783 faktum 154
11784 faktumet 1
11785 falerner 1
11786 fall 283
11787 falla 9
11788 fallen 11
11789 fallenhet 1
11790 faller 24
11791 fallerar 1
11792 fallet 110
11793 fallfärdiga 1
11794 fallfärdigt 1
11795 fallit 10
11796 fallna 1
11797 fallstudie 1
11798 falsk 4
11799 falska 12
11800 falskheten 1
11801 falskmyntare 1
11802 falskmyntarna 1
11803 falskmynteri 1
11804 falskmyntning 3
11805 falskt 2
11806 familj 10
11807 familje- 2
11808 familjeansvaret 3
11809 familjeenheten 1
11810 familjefader 1
11811 familjeförhållandena 1
11812 familjeförändringar 1
11813 familjejordbruk 3
11814 familjejordbruken 1
11815 familjeliv 1
11816 familjelivet 1
11817 familjemedlem 1
11818 familjen 18
11819 familjens 1
11820 familjeovänliga 1
11821 familjepolitik 2
11822 familjer 25
11823 familjerna 1
11824 familjernas 1
11825 familjeägodelar 1
11826 familjeåterförening 2
11827 famn 2
11828 famnen 3
11829 fanan 1
11830 fanatisk 1
11831 fanatiska 1
11832 fann 12
11833 fanns 113
11834 fansen 1
11835 fanstyg 1
11836 fantasi 4
11837 fantasibilder 1
11838 fantasier 1
11839 fantasifulla 2
11840 fantasilösa 1
11841 fantasin 3
11842 fantasirik 1
11843 fantastisk 4
11844 fantastiska 10
11845 fantastiskt 7
11846 fantom 1
11847 fanér 1
11848 far 53
11849 fara 28
11850 faran 6
11851 farbar 1
11852 farbror 4
11853 farfarsfars 1
11854 farföräldrar 2
11855 farföräldrars 1
11856 farhågor 10
11857 farkost 2
11858 farkosten 1
11859 farleden 1
11860 farlig 12
11861 farliga 39
11862 farligare 1
11863 farligaste 1
11864 farligheterna 1
11865 farligt 53
11866 farmakologiska 1
11867 farmor 24
11868 farmors 3
11869 farofyllda 1
11870 faror 5
11871 farorna 2
11872 farozon 1
11873 fars 7
11874 farsartade 1
11875 farsot 1
11876 farsoten 1
11877 farsoter 1
11878 fart 8
11879 farten 1
11880 fartyg 62
11881 fartygen 23
11882 fartygens 8
11883 fartyget 18
11884 fartygets 3
11885 fartygs 3
11886 fartygsavfall 1
11887 fartygsbesättningar 1
11888 fartygsgenererade 1
11889 fartygsgenererat 4
11890 fartygsinspektionen 1
11891 fartygsinspektionsbolaget 1
11892 fartygsolyckan 2
11893 fartygsolyckor 1
11894 fartygssidorna 1
11895 fartygsskrov 9
11896 fartygssäkerhet 2
11897 fartygssäkerheten 1
11898 fartygstankrarna 1
11899 fartygsägaren 1
11900 farvatten 14
11901 fas 15
11902 fasa 2
11903 fasaden 1
11904 fasansfull 1
11905 fasansfulla 2
11906 fasat 1
11907 fascinerade 1
11908 fascineras 1
11909 fascism 2
11910 fascismen 1
11911 fascismens 1
11912 fascistdiktators 1
11913 fascisterna 2
11914 fascisternas 1
11915 fascistisk 1
11916 fascistiska 1
11917 fascistiskt 2
11918 fasen 4
11919 faser 2
11920 faserna 2
11921 fasor 1
11922 fast 97
11923 fasta 18
11924 fasthet 2
11925 fastigheten 1
11926 fastklamrade 1
11927 fastklängda 1
11928 fastkubikmeter 1
11929 fastlagd 1
11930 fastlagda 1
11931 fastlagt 1
11932 fastlagts 2
11933 fastland 2
11934 fastlandet 5
11935 fastlägga 1
11936 fastläggas 1
11937 fastläggs 1
11938 fastnade 1
11939 fastnar 2
11940 fastnat 2
11941 fastsatt 1
11942 fastslagen 1
11943 fastslaget 1
11944 fastslagit 1
11945 fastslagits 2
11946 fastslagna 1
11947 fastslog 4
11948 fastslogs 2
11949 fastslå 9
11950 fastslår 6
11951 fastslås 14
11952 fastställa 60
11953 fastställande 13
11954 fastställandet 4
11955 fastställas 9
11956 fastställd 4
11957 fastställda 8
11958 fastställde 3
11959 fastställdes 10
11960 fastställer 17
11961 fastställs 19
11962 fastställt 6
11963 fastställts 17
11964 fastän 7
11965 fatala 1
11966 fatalitet 1
11967 fatalt 2
11968 fatet 1
11969 fatt 1
11970 fatta 54
11971 fattade 14
11972 fattades 9
11973 fattar 16
11974 fattas 32
11975 fattat 4
11976 fattats 14
11977 fattig 1
11978 fattiga 42
11979 fattigare 6
11980 fattigaste 19
11981 fattigbasaren 2
11982 fattigdom 36
11983 fattigdomen 30
11984 fattigdomsbekämpning 1
11985 fattigdomsbekämpningen 1
11986 fattigdomsbekämpningens 1
11987 fattigdomsdrabbade 1
11988 fattigdomsfokusering 1
11989 fattigdomsgräns 1
11990 fattigdomsgränsen 1
11991 fattigdomsgränser 2
11992 fattigdomsproblematiken 1
11993 fattigdomsproblemen 1
11994 fattigmat 1
11995 fattigt 1
11996 fattning 1
11997 fauna 2
11998 favelas 1
11999 favoritlektyr 1
12000 favör 1
12001 fax 2
12002 faxa 1
12003 fe 1
12004 feber 1
12005 febrigt 1
12006 februari 49
12007 fedayeens 1
12008 federal 6
12009 federala 3
12010 federalism 4
12011 federalist 1
12012 federalister 1
12013 federalisterna 1
12014 federalistisk 3
12015 federalistiska 2
12016 federalt 3
12017 federation 3
12018 federationen 2
12019 federationens 1
12020 federationskärna 1
12021 fee 1
12022 fee-system 1
12023 fee-systemet 2
12024 fel 56
12025 felaktig 9
12026 felaktiga 2
12027 felaktigare 1
12028 felaktighet 1
12029 felaktigheter 2
12030 felaktigt 21
12031 felande 1
12032 felar 1
12033 felberäkning 1
12034 felciterad 1
12035 felet 1
12036 felfritt 1
12037 felkvot 1
12038 felringning 1
12039 felräkningen 1
12040 felsyn 1
12041 feltolkat 1
12042 felöversättning 2
12043 fem 101
12044 femdubblats 1
12045 femfaldigat 1
12046 femminuterssändning 1
12047 fempunktsprogram 1
12048 femte 21
12049 femtedel 3
12050 femtedelar 1
12051 femtedelen 1
12052 femti 1
12053 femtielfte 1
12054 femtio 10
12055 femtioelfte 1
12056 femtioelva 1
12057 femtiotal 1
12058 femtioårsperiodens 1
12059 femton 37
12060 femtonhundra 1
12061 femtonhundratalet 1
12062 femåriga 1
12063 femårigt 1
12064 femårsperiod 7
12065 femårsperioden 1
12066 femårsplan 2
12067 femårsplanen 5
12068 femårsplaner 2
12069 femårsprogram 8
12070 femårsprogrammet 3
12071 fenomen 13
12072 fenomenet 4
12073 fernissade 1
12074 fest 5
12075 fester 1
12076 festerna 2
12077 festkvällar 1
12078 festligheterna 3
12079 festligt 1
12080 festregeln 1
12081 feststämning 1
12082 fet 2
12083 feta 4
12084 fetade 1
12085 fiaskona 1
12086 fiaskot 1
12087 fick 158
12088 ficka 1
12089 fickan 6
12090 fickor 1
12091 fickorna 3
12092 fiducia 1
12093 fiende 5
12094 fiender 6
12095 fiendishly 1
12096 fiendskap 1
12097 fientlig 1
12098 fientliga 3
12099 fientligheterna 3
12100 fientligt 1
12101 figur 1
12102 fikar 1
12103 fil 4
12104 filantropi 1
12105 filen 7
12106 filer 4
12107 filerna 1
12108 filformat 2
12109 filformatet 1
12110 film 1
12111 filmdukar 1
12112 filmen 1
12113 filmens 1
12114 filmer 1
12115 filmerna 1
12116 filmsuccé 1
12117 filoberoende 1
12118 filosof 1
12119 filosofi 9
12120 filosofibok 1
12121 filosofin 2
12122 filosofisk 2
12123 filosofiska 2
12124 filtar 3
12125 filten 1
12126 filter 14
12127 filteraxeln 1
12128 filterfunktioner 1
12129 filterfält 3
12130 filterfältet 1
12131 filterinställningar 1
12132 filterinställningarna 1
12133 filterområdet 3
12134 filterval 1
12135 filtrera 14
12136 filtrerade 1
12137 filtrerar 4
12138 filtreras 2
12139 filtrerat 2
12140 filtrering 3
12141 filtreringen 2
12142 filtret 3
12143 fin 1
12144 fina 9
12145 finans 1
12146 finans- 1
12147 finansdepartementet 1
12148 finanser 5
12149 finanseringsreformen 1
12150 finanserna 2
12151 finansernas 1
12152 finansföretagens 1
12153 finansgrupp 1
12154 finansiell 12
12155 finansiella 75
12156 finansiellt 17
12157 finansiera 31
12158 finansierad 2
12159 finansierade 3
12160 finansierar 5
12161 finansieras 25
12162 finansierat 2
12163 finansierats 3
12164 finansiering 35
12165 finansieringen 31
12166 finansieringsbeloppet 1
12167 finansieringsbidrag 1
12168 finansieringsinstrument 1
12169 finansieringsinstrumentet 2
12170 finansieringskapital 1
12171 finansieringskällor 1
12172 finansieringsmarknaden 1
12173 finansieringsmetoder 1
12174 finansieringsmodell 1
12175 finansieringsmöjligheter 1
12176 finansieringspaketet 1
12177 finansieringsplan 1
12178 finansieringsplanerna 1
12179 finansieringsprogram 1
12180 finansieringsramar 1
12181 finansieringsramen 1
12182 finansieringsstöd 1
12183 finansieringssystemen 1
12184 finansieringstjänster 1
12185 finansieringsvolym 2
12186 finansieringsåtgärder 1
12187 finansinstituten 2
12188 finansinstrument 1
12189 finansiärer 2
12190 finansiärerna 2
12191 finansmarknaderna 1
12192 finansmarknadernas 1
12193 finansmedlen 1
12194 finansminister 2
12195 finansministern 4
12196 finansministerns 1
12197 finansministrarna 1
12198 finansmän 1
12199 finanspolitik 1
12200 finansprogram 1
12201 finansprotokoll 1
12202 finansprotokollen 2
12203 finansredskap 1
12204 finanssystem 1
12205 finanstekniska 1
12206 finansutskott 1
12207 finaste 2
12208 finding 1
12209 finesse 1
12210 finesser 1
12211 finfördela 1
12212 finge 1
12213 finger 1
12214 fingeravtrycken 1
12215 fingervisning 2
12216 fingrar 3
12217 fingrarna 4
12218 fingret 2
12219 finhet 1
12220 finkänsliga 1
12221 finkänsligt 1
12222 finländare 1
12223 finländska 9
12224 finn 1
12225 finna 58
12226 finnar 1
12227 finnas 112
12228 finner 28
12229 finnig 1
12230 finns 944
12231 finsk 4
12232 finska 10
12233 finskuren 1
12234 finskurna 1
12235 fint 2
12236 fira 4
12237 firade 1
12238 firandet 2
12239 firma 1
12240 firman 2
12241 fisk 26
12242 fiska 12
12243 fiskades 1
12244 fiskar 11
12245 fiskare 12
12246 fiskaren 2
12247 fiskarna 11
12248 fiskarnas 2
12249 fiskarter 5
12250 fiskas 1
12251 fiskats 1
12252 fiskbankar 1
12253 fiskbestånd 5
12254 fiskbestånden 5
12255 fiskbeståndet 2
12256 fiske 36
12257 fiske- 3
12258 fiskeansträngningar 1
12259 fiskeansträngningarna 1
12260 fiskeansträngningen 1
12261 fiskeavtalen 1
12262 fiskebankarna 1
12263 fiskeby 1
12264 fiskebåtar 1
12265 fiskedagarna 1
12266 fiskefartyg 3
12267 fiskefartyget 1
12268 fiskeflotta 2
12269 fiskeflottan 1
12270 fiskeflottor 1
12271 fiskefrågan 1
12272 fiskeindustrins 1
12273 fiskekvoterna 1
12274 fiskelivet 1
12275 fiskemetodernas 1
12276 fiskemängden 1
12277 fiskemöjligheter 4
12278 fisken 8
12279 fiskens 1
12280 fiskeodlingar 1
12281 fiskeområde 1
12282 fiskeområdet 1
12283 fiskeorganisationerna 1
12284 fiskepolitik 1
12285 fiskeprodukter 1
12286 fiskeprodukterna 1
12287 fiskeproduktionen 2
12288 fiskeredskap 2
12289 fiskeredskapen 2
12290 fiskeregion 1
12291 fiskeresurser 1
12292 fiskeresurserna 10
12293 fiskeriansträngningarna 1
12294 fiskeriet 3
12295 fiskerifrågor 1
12296 fiskeriförvaltning 3
12297 fiskeriindustri 1
12298 fiskeriindustrin 1
12299 fiskerikommittén 1
12300 fiskerilagstiftningen 1
12301 fiskerinäring 1
12302 fiskerinäringen 9
12303 fiskerinäringens 1
12304 fiskeriområdet 3
12305 fiskeriorganisation 1
12306 fiskeriorganisationerna 4
12307 fiskeripolitik 10
12308 fiskeripolitiken 35
12309 fiskeripolitikens 2
12310 fiskeriresurserna 1
12311 fiskerisektor 3
12312 fiskerisektorer 1
12313 fiskerisektorn 23
12314 fiskeristatistiken 1
12315 fiskeriutskott 3
12316 fiskeriutskottet 26
12317 fiskeriutskottets 2
12318 fiskeriverksamhet 6
12319 fiskeriverksamheten 6
12320 fiskerättigheter 2
12321 fiskesamhällen 3
12322 fiskesamhällenas 1
12323 fiskesektorer 1
12324 fiskesektorn 4
12325 fiskestopp 1
12326 fisket 39
12327 fisketrycket 3
12328 fiskets 3
12329 fiskeuppgifter 1
12330 fiskevattnen 2
12331 fiskeverksamheten 1
12332 fiskfångst 1
12333 fiskfångstfartyg 1
12334 fiskgrossister 1
12335 fiskodling 3
12336 fiskodlingar 1
12337 fiskodlingen 1
12338 fiskodlingssektorn 1
12339 fiskprodukter 1
12340 fisksjukdomar 2
12341 fission 1
12342 fixa 1
12343 fixera 1
12344 fjol 6
12345 fjolårets 1
12346 fjorton 17
12347 fjortonde 1
12348 fjortonsidiga 1
12349 fjädrarna 1
12350 fjärde 37
12351 fjärde- 1
12352 fjärdedel 3
12353 fjärdedelar 3
12354 fjärilarna 1
12355 fjärma 1
12356 fjärmade 1
12357 fjärran 2
12358 flacka 1
12359 fladdermusliknande 1
12360 fladdrande 2
12361 flagg 10
12362 flagga 5
12363 flaggan 2
12364 flaggens 1
12365 flaggorna 1
12366 flaggskepp 1
12367 flaggstång 1
12368 flagnande 1
12369 flagrant 2
12370 flamländska 2
12371 flammade 1
12372 flammat 1
12373 flammorna 1
12374 flampulver 2
12375 flamskyddsmedel 5
12376 flamskyddsmedlen 1
12377 flaska 5
12378 flaskan 3
12379 flaskhals 1
12380 flaskor 2
12381 flaskorna 1
12382 flaxade 1
12383 fleece 1
12384 fler 77
12385 flera 224
12386 flerstatlig 1
12387 flertal 12
12388 flertalet 11
12389 flerårig 3
12390 fleråriga 9
12391 flerårigt 8
12392 flerårsbasis 1
12393 flerårsbudget 1
12394 flesta 60
12395 flexibel 15
12396 flexibelt 13
12397 flexibilisering 1
12398 flexibilitet 36
12399 flexibiliteten 3
12400 flexibilitetsklausul 2
12401 flexibla 12
12402 flexiblare 3
12403 flexible 1
12404 flicka 7
12405 flickan 6
12406 flickans 1
12407 flickor 6
12408 flickorna 3
12409 flickors 1
12410 flimmer 1
12411 flimret 1
12412 flin 1
12413 flinade 2
12414 flingor 2
12415 flintskallig 2
12416 flirta 1
12417 flit 2
12418 fliten 1
12419 flitigare 1
12420 flock 1
12421 flod 7
12422 flod-team 1
12423 flodarm 1
12424 flodbåt 1
12425 floden 29
12426 flodens 1
12427 floder 8
12428 floderna 3
12429 flodernas 2
12430 floders 1
12431 flodledens 1
12432 flodmynningen 3
12433 flodstränder 1
12434 flodstränderna 1
12435 flodvattendistrikt 1
12436 flodvattendistrikten 1
12437 flodvattnet 1
12438 flodvåg 1
12439 flora 2
12440 florida 1
12441 flottan 5
12442 flottans 1
12443 flottiga 1
12444 flottigt 1
12445 flottkapacitet 1
12446 flottkapaciteten 1
12447 flottorna 2
12448 fluff 1
12449 fluga 1
12450 flugit 1
12451 flugor 3
12452 fluktuationsmarginal 1
12453 flutit 1
12454 fly 2
12455 flydde 3
12456 flyg 6
12457 flyga 6
12458 flygande 4
12459 flyganfall 1
12460 flygbiljett 1
12461 flygblad 1
12462 flygbolag 2
12463 flygbombningarna 1
12464 flyger 2
12465 flyget 3
12466 flygkrascherna 1
12467 flyglinjerna 1
12468 flygningen 1
12469 flygplan 3
12470 flygplanen 1
12471 flygplanet 1
12472 flygplanskerosin 1
12473 flygplats 2
12474 flygplatsen 4
12475 flygplatser 2
12476 flygpriserna 1
12477 flygräd 1
12478 flygs 1
12479 flygsäkerheten 1
12480 flygtransport 1
12481 flygtransporter 2
12482 flygtransporterna 1
12483 flygturer 1
12484 flygvärdinnan 1
12485 flykt 5
12486 flykten 5
12487 flyktig 1
12488 flykting 2
12489 flykting- 1
12490 flyktingar 30
12491 flyktingarna 8
12492 flyktingeländet 1
12493 flyktingfonden 1
12494 flyktingfrågor 1
12495 flyktingkommissariat 2
12496 flyktingpolitik 3
12497 flyktingpolitiken 2
12498 flyktingskollärare 1
12499 flyktingstatus 5
12500 flyktingströmmarnas 1
12501 flyktingstödet 1
12502 flyktmöjlighet 1
12503 flyr 1
12504 flyta 1
12505 flytande 1
12506 flyter 2
12507 flytet 1
12508 flytetyg 1
12509 flytt 3
12510 flytta 29
12511 flyttade 9
12512 flyttar 16
12513 flyttas 12
12514 flyttat 5
12515 flyttats 1
12516 flyttfåglar 1
12517 flyttningen 1
12518 flyttningsprogram 1
12519 flyttningsprogrammet 1
12520 fläck 5
12521 fläckar 3
12522 fläcken 2
12523 fläckigt 1
12524 fläkt 2
12525 fläktarna 2
12526 flämtade 3
12527 flämtande 2
12528 fläng 1
12529 flå 1
12530 flåsande 4
12531 flöde 1
12532 flöden 2
12533 flödet 3
12534 flödiga 1
12535 flög 7
12536 flöjt 1
12537 flörtade 1
12538 flörtig 1
12539 flöt 5
12540 foder 10
12541 foderantibiotika 1
12542 foderblandningar 2
12543 foderdirektivet 1
12544 fodermaterial 1
12545 fodertillsatsen 1
12546 fodertillsatser 14
12547 fodertillsatserna 3
12548 fodertillverkares 1
12549 fog 1
12550 foga 2
12551 fogades 1
12552 fogas 1
12553 fogat 3
12554 foie 3
12555 fokus 5
12556 fokusera 7
12557 fokuserar 7
12558 fokuseras 2
12559 fokuserat 1
12560 fokusering 5
12561 fokuseringen 1
12562 folk 74
12563 folkbibliotek 1
12564 folken 8
12565 folkens 9
12566 folket 27
12567 folketing 1
12568 folketinget 2
12569 folkets 13
12570 folkgrupp 1
12571 folkgrupper 2
12572 folkgrupperna 7
12573 folkhälsa 29
12574 folkhälsan 13
12575 folkhälsans 1
12576 folkhälsoaspekterna 1
12577 folkhälsofråga 2
12578 folkhälsoplanet 1
12579 folkhälsorisk 1
12580 folkhälsoskäl 1
12581 folklagren 2
12582 folklore 1
12583 folkmassan 4
12584 folkmord 7
12585 folkmyllret 2
12586 folkomröstning 5
12587 folkomröstningar 3
12588 folkomröstningen 1
12589 folkopinion 1
12590 folkpartiet 16
12591 folkpartiets 26
12592 folkregeringar 1
12593 folkrepublikens 1
12594 folkräkning 1
12595 folkräkningen 1
12596 folkrätt 1
12597 folkrätten 3
12598 folkrörelserna 1
12599 folks 7
12600 folkskolorna 1
12601 folkstyrets 1
12602 folksägner 1
12603 folktomt 1
12604 folkvalda 12
12605 folkvaldas 1
12606 fond 12
12607 fondandelar 1
12608 fondbolagen 1
12609 fonden 8
12610 fonder 32
12611 fonderna 15
12612 fondernas 1
12613 fondföretag 14
12614 fondföretagen 6
12615 fondföretagens 2
12616 fondföretagsinvesteringar 1
12617 fondförvaltare 2
12618 fondmedel 3
12619 fonduppbyggnad 1
12620 foots 1
12621 for 15
12622 fora 3
12623 force 3
12624 forcerade 1
12625 fordon 61
12626 fordonen 8
12627 fordonet 2
12628 fordons 1
12629 fordonsindustrin 1
12630 fordonsmärken 1
12631 fordonspark 1
12632 fordonstillverkare 1
12633 fordonstillverkarna 2
12634 fordonsägaren 1
12635 fordonsåtervinningen 1
12636 fordra 1
12637 fordrande 1
12638 fordrar 3
12639 fordras 10
12640 fordringar 1
12641 forell 2
12642 form 104
12643 forma 1
12644 formad 1
12645 formalism 1
12646 formalitet 3
12647 formaliteter 2
12648 formandet 1
12649 formar 1
12650 format 10
12651 formatera 1
12652 formatering 2
12653 formateringen 3
12654 formationer 1
12655 formatmall 1
12656 formatmallar 1
12657 formats 2
12658 formel 3
12659 formell 9
12660 formella 6
12661 formellt 21
12662 formen 8
12663 former 35
12664 formering 1
12665 formerna 6
12666 formulera 10
12667 formulerad 1
12668 formulerade 8
12669 formulerades 2
12670 formuleras 7
12671 formulerat 3
12672 formulerats 6
12673 formulering 7
12674 formuleringar 5
12675 formuleringarna 1
12676 formuleringen 6
12677 formulär 21
12678 formuläret 1
12679 formulärets 2
12680 forna 3
12681 fornminnena 1
12682 forsar 1
12683 forsarna 1
12684 forska 1
12685 forskare 8
12686 forskares 1
12687 forskning 72
12688 forskningen 9
12689 forskningens 2
12690 forsknings- 2
12691 forskningsaktiviteterna 1
12692 forskningsarbeten 1
12693 forskningsbidrag 1
12694 forskningsinformation 1
12695 forskningsinfrastrukturen 1
12696 forskningsområde 4
12697 forskningsområdet 1
12698 forskningsplats 1
12699 forskningspolitik 2
12700 forskningsprogram 5
12701 forskningsprogrammen 1
12702 fort 20
12703 fortare 1
12704 fortbildning 10
12705 fortbildningsprogram 1
12706 fortet 1
12707 fortfarande 307
12708 fortgå 7
12709 fortgående 6
12710 fortlevnad 2
12711 fortlöpande 5
12712 fortlöper 1
12713 fortplantas 1
12714 fortsatt 21
12715 fortsatta 12
12716 fortsatte 18
12717 fortskaffningsmedel 1
12718 fortskrida 1
12719 fortskridande 2
12720 fortskrider 3
12721 fortsätt 2
12722 fortsätta 135
12723 fortsättas 1
12724 fortsätter 82
12725 fortsättning 15
12726 fortsättningen 28
12727 fortsättningsvis 4
12728 forum 8
12729 forumet 5
12730 forêts 1
12731 fosfor 1
12732 fosforrött 1
12733 fossila 2
12734 fosterland 2
12735 fot 7
12736 fotboll 1
12737 fotbollsbedrägerierna 1
12738 fotbollsplan 1
12739 foten 4
12740 fotfäste 1
12741 fotgängarna 1
12742 fotoförstoringar 1
12743 fotograferade 1
12744 fotografi 6
12745 fotografier 2
12746 fotografiet 2
12747 fotona 1
12748 fotot 1
12749 fots 2
12750 fotspår 2
12751 fotsvamp 1
12752 fotvärmare 1
12753 frack 1
12754 fragment 1
12755 fragmentariskt 1
12756 fragmenterade 1
12757 frakta 1
12758 fraktats 1
12759 fraktens 2
12760 fraktfartyg 1
12761 fraktfordon 1
12762 fram 706
12763 frambesvärja 1
12764 frambringade 1
12765 frambringar 1
12766 framdeles 5
12767 framfart 2
12768 framfusigt 1
12769 framfödde 1
12770 framför 325
12771 framföra 42
12772 framförallt 1
12773 framförande 1
12774 framföranden 3
12775 framföras 1
12776 framförd 1
12777 framförde 13
12778 framförhandlad 1
12779 framförhandlas 1
12780 framförhandlats 1
12781 framförs 7
12782 framfört 12
12783 framförts 17
12784 framgick 4
12785 framgå 3
12786 framgång 47
12787 framgångar 13
12788 framgångarna 2
12789 framgångarnas 1
12790 framgången 7
12791 framgångens 1
12792 framgångsfaktor 1
12793 framgångsrik 19
12794 framgångsrika 12
12795 framgångsrikt 19
12796 framgångssagor 1
12797 framgår 26
12798 framgått 2
12799 framhärda 1
12800 framhärdandet 1
12801 framhärdar 1
12802 framhäva 4
12803 framhävas 2
12804 framhävde 1
12805 framhäver 1
12806 framhävs 2
12807 framhävt 1
12808 framhålla 25
12809 framhållas 2
12810 framhåller 12
12811 framhållit 8
12812 framhålls 2
12813 framhöll 6
12814 framhölls 1
12815 framkalla 2
12816 framkallade 2
12817 framkallar 1
12818 framkallat 5
12819 framkastat 1
12820 framkom 3
12821 framkommer 8
12822 framkommit 7
12823 framlade 1
12824 framlagda 8
12825 framlagt 5
12826 framlagts 6
12827 framlägga 2
12828 framläggandet 3
12829 framlägger 2
12830 framläggs 2
12831 frammana 1
12832 framme 3
12833 framröstade 1
12834 framsida 1
12835 framsidan 1
12836 framskjuten 1
12837 framskjutna 2
12838 framskrider 1
12839 framskridet 1
12840 framskridna 1
12841 framsteg 86
12842 framstegen 7
12843 framsteget 2
12844 framstod 1
12845 framställa 9
12846 framställan 1
12847 framställd 1
12848 framställde 1
12849 framställer 1
12850 framställning 10
12851 framställningar 9
12852 framställningarna 1
12853 framställningen 2
12854 framställs 3
12855 framställt 1
12856 framställts 2
12857 framstå 2
12858 framstående 10
12859 framstår 6
12860 framstötar 1
12861 framsätet 2
12862 framtagandet 4
12863 framtagits 1
12864 framtagning 1
12865 framtid 60
12866 framtida 63
12867 framtiden 148
12868 framtidens 4
12869 framtidsbild 1
12870 framtidsdugliga 1
12871 framtidsförmåga 1
12872 framtidshopp 1
12873 framtidsinriktad 1
12874 framtidsinriktat 1
12875 framtidsorienterad 1
12876 framtidsorienterat 1
12877 framtidsutsikter 5
12878 framtidsutsikterna 1
12879 framtoning 1
12880 framträda 2
12881 framträdande 7
12882 framträder 5
12883 framtvingade 1
12884 framtvingar 1
12885 framtvingas 2
12886 framtvingbara 1
12887 framväxande 3
12888 framväxten 1
12889 framåt 66
12890 framåtböjd 1
12891 framåtmarsch 1
12892 framåtskridande 1
12893 framöver 12
12894 franc 5
12895 franca 1
12896 franchisesystem 1
12897 frankiskt 1
12898 fransk 5
12899 franska 76
12900 franske 3
12901 franskt 2
12902 fransktalande 1
12903 franskägt 1
12904 fransmän 1
12905 fransmännen 5
12906 frapperande 1
12907 fras 1
12908 frasen 1
12909 fraser 1
12910 frasig 1
12911 fred 66
12912 fredag 7
12913 fredagen 3
12914 freden 20
12915 fredens 4
12916 fredlig 13
12917 fredliga 4
12918 fredligt 4
12919 fredsansträngningar 1
12920 fredsavtal 6
12921 fredsavtalen 1
12922 fredsavtalet 4
12923 fredsbeskyddare 1
12924 fredsbevarande 6
12925 fredsbyggande 2
12926 fredsbyggare 1
12927 fredsfrämjande 1
12928 fredsförhandlingarna 3
12929 fredsgrupper 1
12930 fredslösning 1
12931 fredsordning 1
12932 fredsorganisationer 1
12933 fredspartner 1
12934 fredsplan 1
12935 fredsprocess 6
12936 fredsprocessen 37
12937 fredsprocessens 2
12938 fredsprocesser 1
12939 fredsrörelse 1
12940 fredssamarbete 1
12941 fredssamtal 1
12942 fredssamtalen 4
12943 fredssituation 1
12944 fredsskapande 1
12945 fredsstiftande 1
12946 fredsstyrka 1
12947 fredsuppgörelse 3
12948 free 1
12949 frekventera 2
12950 frenetiskt 1
12951 fresker 1
12952 fresta 1
12953 frestas 1
12954 frestelsen 3
12955 fri 47
12956 fri- 32
12957 fria 68
12958 friare 1
12959 friat 1
12960 frid 4
12961 friden 1
12962 fridfullt 1
12963 fridsamt 1
12964 frigiven 1
12965 frigivningen 1
12966 frigjorda 1
12967 frigjordhet 1
12968 frigjort 1
12969 frigör 1
12970 frigöra 8
12971 frigörande 1
12972 frigöras 1
12973 frigörs 1
12974 frihandel 1
12975 frihandeln 1
12976 frihandelns 4
12977 frihandelsavtalen 1
12978 frihandelsområde 1
12979 frihandelsområden 1
12980 frihandelsområdena 1
12981 frihandelspolitiken 1
12982 frihandelsuppgörelser 1
12983 frihandelsvänliga 1
12984 frihandelszon 1
12985 frihet 97
12986 friheten 20
12987 frihetens 5
12988 friheter 11
12989 friheterna 8
12990 frihetsberövad 1
12991 frihetsberövande 1
12992 frihetskamp 1
12993 frihetskänsla 1
12994 frihetsparti 1
12995 frikostigt 2
12996 friktionsfria 1
12997 frilansande 1
12998 frimurarna 2
12999 frimärken 1
13000 frimärkspriser 1
13001 frisersalong 1
13002 frisk 3
13003 friska 3
13004 friskt 2
13005 frisläppande 3
13006 frisläppandet 1
13007 frisläppt 1
13008 fristaten 1
13009 fristen 1
13010 frister 2
13011 friställningar 1
13012 fristående 3
13013 frisördockas 1
13014 fritid 1
13015 fritids- 1
13016 fritidssituationer 1
13017 fritidssysselsättningar 1
13018 fritt 18
13019 frivillig 5
13020 frivillig- 1
13021 frivilliga 14
13022 frivilligas 1
13023 frivilligorganisationer 1
13024 frivilligsektorn 1
13025 frivilligt 7
13026 frodas 6
13027 from 1
13028 fromhet 1
13029 fromma 3
13030 front 1
13031 frontalangreppet 1
13032 fronten 4
13033 fronter 1
13034 frontlinjen 1
13035 frost 1
13036 frosten 1
13037 fru 169
13038 fruar 1
13039 frukost 4
13040 frukostbordet 1
13041 frukosten 2
13042 frukostägg 1
13043 frukt 4
13044 fruktade 3
13045 fruktades 1
13046 fruktan 5
13047 fruktande 1
13048 fruktansvärd 5
13049 fruktansvärda 10
13050 fruktansvärt 6
13051 fruktar 13
13052 fruktat 1
13053 fruktbara 1
13054 fruktbart 7
13055 fruktbiffar 1
13056 frukten 3
13057 fruktkaka 1
13058 fruktsamhet 1
13059 fruntimmer 1
13060 frusenheten 1
13061 frusna 1
13062 frustade 1
13063 frustar 2
13064 frustration 4
13065 frustrationen 2
13066 frustrerade 1
13067 frustrering 1
13068 frysa 2
13069 frysen 1
13070 fräckhet 1
13071 fräckheten 1
13072 fräkniga 1
13073 fräknigt 1
13074 främja 117
13075 främjade 2
13076 främjande 16
13077 främjandet 11
13078 främjar 32
13079 främjare 1
13080 främjas 8
13081 främjat 3
13082 främling 2
13083 främlingar 3
13084 främlingen 2
13085 främlingens 1
13086 främlings- 1
13087 främlingsfientlig 2
13088 främlingsfientliga 23
13089 främlingsfientlighet 25
13090 främlingsfientligheten 2
13091 främlingsfientlighetens 2
13092 främlingsfientligt 5
13093 främlingshat 1
13094 främlingsrädsla 1
13095 främlingsskap 1
13096 främmande 13
13097 främst 97
13098 främsta 39
13099 främste 2
13100 fräsanden 1
13101 fräsch 1
13102 fräste 1
13103 fråga 789
13104 frågade 31
13105 frågan 489
13106 frågande 6
13107 frågans 4
13108 frågar 51
13109 frågat 6
13110 frågekomplex 1
13111 frågeläge 5
13112 frågelägen 1
13113 frågelägesinställning 1
13114 frågeläget 1
13115 frågesatsen 1
13116 frågestunden 15
13117 frågeställaren 4
13118 frågeställningen 1
13119 frågetecken 4
13120 frågor 496
13121 frågorna 74
13122 från 1917
13123 frångår 1
13124 frånsett 1
13125 frånstötande 1
13126 frånsäga 1
13127 fråntar 1
13128 fråntas 3
13129 fråntog 1
13130 frånvarande 15
13131 frånvaro 8
13132 frånvaron 6
13133 frö 2
13134 fröet 1
13135 fröjdar 1
13136 fukt 1
13137 fuktigt 1
13138 fulhet 1
13139 full 76
13140 fulla 25
13141 fullare 1
13142 fullaste 1
13143 fullborda 3
13144 fullbordad 3
13145 fullbordandet 2
13146 fullbordar 1
13147 fullbordas 2
13148 fullbordat 1
13149 fullfölja 4
13150 fullföljas 1
13151 fullföljer 3
13152 fullföljt 1
13153 fullgjort 2
13154 fullgör 1
13155 fullgöra 7
13156 fullgöras 2
13157 fullgörs 1
13158 fullkomlig 1
13159 fullkomlighet 1
13160 fullkomligt 9
13161 fullkomnade 1
13162 fullmakt 2
13163 fullmaktsbestämmelser 1
13164 fullmäktige 1
13165 fullo 8
13166 fullpackad 1
13167 fullsatt 1
13168 fullständig 34
13169 fullständiga 11
13170 fullständigt 71
13171 fullt 62
13172 fulltecknade 1
13173 fulltoniga 1
13174 fullvärdig 6
13175 fullvärdiga 2
13176 fullända 1
13177 fulländar 1
13178 fulländat 1
13179 fult 1
13180 fumlig 1
13181 fundamental 1
13182 fundamentala 2
13183 fundamentalt 3
13184 fundera 18
13185 funderade 9
13186 funderar 8
13187 funderingar 3
13188 funderingarna 1
13189 fundersökningar 1
13190 fungera 56
13191 fungerade 3
13192 fungerande 23
13193 fungerar 59
13194 fungerat 8
13195 funktion 31
13196 funktionalistiska 2
13197 funktionella 1
13198 funktionellt 1
13199 funktionen 7
13200 funktioner 13
13201 funktionerna 4
13202 funktionsbrister 1
13203 funktionsduglig 1
13204 funktionsduglighet 3
13205 funktionshinder 8
13206 funktionsregler 2
13207 funktionssätt 1
13208 funktionsvillkor 1
13209 funktionärer 1
13210 funktionärers 1
13211 funnit 9
13212 funnits 24
13213 fusion 2
13214 fusionen 2
13215 fusioner 9
13216 fusionsförordningen 1
13217 fusionshaussen 1
13218 fusionskontrollen 1
13219 fusionsrätten 1
13220 fusk 1
13221 futtiga 2
13222 fylla 14
13223 fyllande 1
13224 fyllas 3
13225 fylld 3
13226 fyllda 2
13227 fyllde 6
13228 fylldes 2
13229 fyller 2
13230 fyllig 2
13231 fylls 1
13232 fyllt 7
13233 fyllts 2
13234 fyra 90
13235 fyrahundra 3
13236 fyratusen 1
13237 fyrkant 1
13238 fyrtio 8
13239 fyrtioett 1
13240 fyrtiosju 1
13241 fyrtiotalet 1
13242 fyrtioåtta 1
13243 fysiken 1
13244 fysiologiska 1
13245 fysisk 9
13246 fysiska 17
13247 fysiskt 7
13248 fädernearvet 1
13249 fällan 1
13250 fällde 2
13251 fäller 1
13252 fälls 1
13253 fällt 1
13254 fällts 3
13255 fält 44
13256 fältelement 1
13257 fälten 7
13258 fältet 27
13259 fältets 2
13260 fängelse 9
13261 fängelsedagbok 1
13262 fängelser 1
13263 fängelserna 3
13264 fängelsestraff 2
13265 fängslas 1
13266 fängslats 1
13267 färd 9
13268 färdades 1
13269 färdats 1
13270 färden 2
13271 färdig 4
13272 färdiga 2
13273 färdigheter 1
13274 färdigställa 1
13275 färdigställde 1
13276 färdigt 8
13277 färdriktning 1
13278 färg 5
13279 färgad 2
13280 färgade 2
13281 färgas 1
13282 färgen 5
13283 färger 8
13284 färgkombinationen 1
13285 färgkänsla 1
13286 färgskrubben 1
13287 färje- 1
13288 färjetrafiken 1
13289 färre 10
13290 färska 1
13291 färskt 2
13292 färskvatten 2
13293 färskvattenförsörjning 1
13294 fäst 4
13295 fästa 9
13296 fästad 1
13297 fästade 1
13298 fäste 1
13299 fäster 8
13300 fästingar 1
13301 fästning 1
13302 fästs 1
13303 få 664
13304 fåfänga 3
13305 fågel 3
13306 fågeldirektiven 1
13307 fågeldirektivet 1
13308 fågellivet 1
13309 fågelpopulationer 1
13310 fågelskrämma 1
13311 fågelskyddssällskapet 1
13312 fågelvänner 1
13313 fåglar 13
13314 fålla 1
13315 fån 1
13316 fånga 1
13317 fångade 4
13318 fångades 1
13319 fångande 1
13320 fångar 13
13321 fångarna 6
13322 fångarnas 1
13323 fångars 1
13324 fångas 1
13325 fångat 3
13326 fånge 1
13327 fångna 2
13328 fångst 5
13329 fångsten 1
13330 fångster 2
13331 fångsterna 2
13332 fångstförbud 1
13333 fångstkvoter 1
13334 fångstmetoder 1
13335 fångstmängd 2
13336 fångstmängden 3
13337 får 582
13338 fårad 1
13339 fåret 1
13340 fårköttsproduktion 1
13341 fåror 1
13342 fås 2
13343 fåtal 10
13344 fåtalet 1
13345 fåtaliga 1
13346 fått 199
13347 fåtölj 1
13348 fåtöljer 1
13349 fåtöljerna 1
13350 föda 2
13351 födande 3
13352 född 2
13353 födda 3
13354 födde 1
13355 föddes 12
13356 födelse 1
13357 födelseakt 1
13358 födelsebygd 1
13359 födelsedag 1
13360 födelsedagen 1
13361 födelsedagshälsningar 1
13362 födelsedagskalasen 1
13363 födelseort 1
13364 födelsetal 1
13365 föder 4
13366 födoämnen 1
13367 föds 4
13368 födsel 2
13369 födseln 1
13370 föga 6
13371 följa 80
13372 följaktligen 36
13373 följande 114
13374 följas 12
13375 följd 68
13376 följde 17
13377 följden 5
13378 följder 14
13379 följderna 12
13380 följdes 5
13381 följdfråga 1
13382 följdfrågan 1
13383 följdfrågor 1
13384 följdriktig 1
13385 följdskador 1
13386 följdskadorna 1
13387 följdåtgärder 1
13388 följe 3
13389 följer 44
13390 följerätten 1
13391 följs 6
13392 följt 16
13393 följts 4
13394 föll 13
13395 fönster 10
13396 fönsterbrädan 2
13397 fönsterbrädet 1
13398 fönstergallret 1
13399 fönsterkarmar 1
13400 fönsterluckorna 1
13401 fönsterlådor 1
13402 fönsterplats 1
13403 fönsterrutorna 1
13404 fönstren 3
13405 fönstret 16
13406 för 9783
13407 föra 82
13408 förakt 3
13409 föraktar 1
13410 föraktat 1
13411 föraktfull 1
13412 föraktfullt 1
13413 föraktlig 1
13414 förankra 2
13415 förankrad 2
13416 förankrade 5
13417 förankras 1
13418 förankring 1
13419 föranleda 1
13420 föranledde 3
13421 föranleder 3
13422 föranslutningsavtal 1
13423 föranslutningsstrategi 2
13424 föranslutningsstrategin 3
13425 föranslutningsstöd 2
13426 förarbetet 1
13427 förare 2
13428 föraren 1
13429 förargat 1
13430 förargligt 1
13431 förarna 2
13432 föras 18
13433 förband 2
13434 förbannat 2
13435 förbannelse 2
13436 förbarmande 1
13437 förbaskat 1
13438 förbehåll 6
13439 förbehållas 3
13440 förbehållen 1
13441 förbehåller 2
13442 förbehållet 1
13443 förbehållslöst 1
13444 förbereda 21
13445 förberedande 14
13446 förberedandet 2
13447 förberedas 5
13448 förberedd 3
13449 förberedda 3
13450 förberedde 4
13451 förbereddes 1
13452 förberedelse 2
13453 förberedelse- 1
13454 förberedelsearbete 1
13455 förberedelsearbetet 1
13456 förberedelsen 2
13457 förberedelseperiod 1
13458 förberedelser 10
13459 förberedelserna 9
13460 förbereder 13
13461 förbereds 2
13462 förberett 4
13463 förberetts 2
13464 förbi 17
13465 förbifarten 2
13466 förbigå 1
13467 förbigående 10
13468 förbigår 1
13469 förbigås 2
13470 förbiilande 1
13471 förbinda 3
13472 förbindelse 14
13473 förbindelselänk 1
13474 förbindelsen 2
13475 förbindelser 40
13476 förbindelseramar 1
13477 förbindelserna 48
13478 förbindelsestrukturen 1
13479 förbinder 8
13480 förbindligheten 1
13481 förbiseende 2
13482 förbisprunget 1
13483 förbisprungits 1
13484 förbittrat 1
13485 förbittring 1
13486 förbjuda 14
13487 förbjudas 5
13488 förbjuden 2
13489 förbjuder 7
13490 förbjudet 7
13491 förbjudit 2
13492 förbjudna 4
13493 förbjuds 1
13494 förbjöd 1
13495 förbjöds 1
13496 förblev 2
13497 förbli 19
13498 förblir 23
13499 förblivande 1
13500 förblivit 1
13501 förbluffade 1
13502 förbluffande 2
13503 förbrukade 1
13504 förbrukar 1
13505 förbrukaren 1
13506 förbrukat 2
13507 förbrukning 2
13508 förbrukningen 1
13509 förbrukningsnivåer 1
13510 förbryllad 1
13511 förbryllande 1
13512 förbrytare 2
13513 förbrytelser 2
13514 förbrytelserna 1
13515 förbränning 1
13516 förbränningskvoten 1
13517 förbränns 1
13518 förbud 18
13519 förbudet 9
13520 förbudsförbehåll 1
13521 förbudsprincipen 1
13522 förbund 1
13523 förbunden 2
13524 förbundet 3
13525 förbundit 9
13526 förbundna 4
13527 förbundskansler 3
13528 förbundskanslern 1
13529 förbundsländer 1
13530 förbundsländerna 1
13531 förbundsregeringen 1
13532 förbundsrepubliken 1
13533 förbättra 107
13534 förbättrad 12
13535 förbättrade 6
13536 förbättrande 1
13537 förbättrar 12
13538 förbättras 19
13539 förbättrat 2
13540 förbättrats 9
13541 förbättring 31
13542 förbättringar 20
13543 förbättringen 4
13544 förbättringstendens 1
13545 förbättringsåtagande 1
13546 förda 3
13547 förde 16
13548 fördefinierade 2
13549 fördel 22
13550 fördela 3
13551 fördelad 1
13552 fördelade 4
13553 fördelaktigt 1
13554 fördelar 19
13555 fördelarna 7
13556 fördelas 7
13557 fördelat 3
13558 fördelats 1
13559 fördelen 4
13560 fördelning 15
13561 fördelningen 9
13562 fördelningsbegreppet 1
13563 fördelningsinstrument 1
13564 fördelningskriterierna 1
13565 fördelningsnyckel 1
13566 fördelningsnyckeln 1
13567 fördelningspolitik 2
13568 fördelningspolitiken 1
13569 fördes 3
13570 fördjupa 12
13571 fördjupad 4
13572 fördjupar 1
13573 fördjupas 2
13574 fördjupat 4
13575 fördjupning 4
13576 fördjupningen 2
13577 fördomar 2
13578 fördomsfrihet 1
13579 fördomsfullhet 1
13580 fördra 2
13581 fördrag 24
13582 fördragen 51
13583 fördragens 5
13584 fördraget 98
13585 fördragets 14
13586 fördrags 1
13587 fördragsanalfabeter 1
13588 fördragsartiklar 1
13589 fördragsfäst 1
13590 fördragsmässiga 1
13591 fördragsmässigt 1
13592 fördragsorganisationens 1
13593 fördragsreform 1
13594 fördragsreglerna 1
13595 fördragssituation 1
13596 fördragsslutande 2
13597 fördragstexten 1
13598 fördragstexterna 1
13599 fördragsändringar 2
13600 fördragsändringarna 1
13601 fördrev 1
13602 fördrivits 1
13603 fördrivna 1
13604 fördrivning 1
13605 fördröja 1
13606 fördröjas 1
13607 fördröjning 1
13608 fördubbla 4
13609 fördubblade 1
13610 fördubblades 1
13611 fördubblas 1
13612 fördubbling 1
13613 fördunklat 1
13614 fördunklats 1
13615 fördämningar 1
13616 fördärva 3
13617 fördärvad 2
13618 fördärvat 1
13619 fördärvbringande 1
13620 fördärvlig 1
13621 fördöma 18
13622 fördömande 11
13623 fördömanden 2
13624 fördömandet 1
13625 fördömas 1
13626 fördömer 17
13627 fördömt 2
13628 fördömts 1
13629 före 103
13630 före-före 1
13631 förebild 9
13632 förebildsmodellen 1
13633 förebråelse 1
13634 förebråelser 1
13635 förebrående 1
13636 förebrås 2
13637 förebygga 18
13638 förebyggande 40
13639 förebyggandet 6
13640 förebyggas 2
13641 förebygger 1
13642 förebådade 1
13643 föredra 11
13644 föredrag 1
13645 föredragande 79
13646 föredraganden 158
13647 föredragandena 8
13648 föredragandenas 1
13649 föredragandens 25
13650 föredragandes 2
13651 föredragit 4
13652 föredragning 2
13653 föredragningslista 18
13654 föredragningslistan 102
13655 föredragningslistor 1
13656 föredragningslistorna 2
13657 föredrar 9
13658 föredrog 3
13659 föredöme 4
13660 föredömlig 1
13661 föredömliga 2
13662 föredömligt 4
13663 förefalla 1
13664 förefaller 45
13665 föreföll 4
13666 föregick 1
13667 föregiven 1
13668 föregripa 2
13669 föregripande 3
13670 föregriper 1
13671 föregripit 1
13672 föregå 3
13673 föregående 57
13674 föregångare 8
13675 föregångares 1
13676 föregångarna 1
13677 föregår 1
13678 föregås 1
13679 förehavanden 3
13680 förekom 3
13681 förekomma 14
13682 förekommande 10
13683 förekommas 1
13684 förekommer 32
13685 förekommit 13
13686 förekomsten 5
13687 förelegat 1
13688 föreligga 2
13689 föreliggande 18
13690 föreligger 29
13691 föreläsa 2
13692 föreläsning 1
13693 föreläsningen 1
13694 föreläste 1
13695 förelåg 1
13696 föremål 38
13697 föremålen 2
13698 föremålet 1
13699 fören 1
13700 förena 25
13701 förenad 2
13702 förenade 4
13703 förenar 4
13704 förenas 3
13705 förenat 1
13706 förenats 1
13707 förening 7
13708 föreningar 3
13709 föreningarna 1
13710 föreningen 1
13711 förenkla 9
13712 förenklad 1
13713 förenklade 4
13714 förenklande 1
13715 förenklar 3
13716 förenklas 1
13717 förenkling 6
13718 förenlig 4
13719 förenliga 7
13720 förenlighet 1
13721 förenligheten 1
13722 förenligt 4
13723 förenta 3
13724 föresats 1
13725 föresatsen 2
13726 föresatser 9
13727 föresatserna 1
13728 föresatt 1
13729 föresatte 1
13730 föreskrev 1
13731 föreskrift 2
13732 föreskrifter 16
13733 föreskrifterna 2
13734 föreskriva 6
13735 föreskrivande 2
13736 föreskriven 1
13737 föreskriver 19
13738 föreskrivit 1
13739 föreskrivits 3
13740 föreskrivna 1
13741 föreskrivs 12
13742 föreslagen 4
13743 föreslagit 40
13744 föreslagits 20
13745 föreslagna 43
13746 föreslog 18
13747 föreslogs 6
13748 föreslå 48
13749 föreslår 88
13750 föreslås 39
13751 förespegla 1
13752 förespeglar 1
13753 förespråka 6
13754 förespråkar 15
13755 förespråkare 6
13756 förespråkarna 2
13757 förespråkas 1
13758 förespråkat 2
13759 förespråkats 1
13760 föreställa 17
13761 föreställde 2
13762 föreställdes 1
13763 föreställer 5
13764 föreställning 1
13765 föreställningar 4
13766 föreställningar- 1
13767 föreställningen 1
13768 föreställt 2
13769 föreståeligt 1
13770 förestående 12
13771 föreståndare 1
13772 föresätter 1
13773 företa 3
13774 företag 212
13775 företagande 4
13776 företagaranda 9
13777 företagarandan 1
13778 företagare 12
13779 företagaren 2
13780 företagarna 7
13781 företagarorganisationer 1
13782 företagartillfällen 1
13783 företagarvärlden 1
13784 företagen 83
13785 företagens 32
13786 företaget 30
13787 företagets 4
13788 företags 3
13789 företags- 1
13790 företagsamhet 10
13791 företagsamma 1
13792 företagsandan 1
13793 företagsavtal 1
13794 företagsbeskattning 1
13795 företagsbeslutet 1
13796 företagsdemokratisering 1
13797 företagsekonomisk 1
13798 företagsekonomiska 3
13799 företagsekonomiskt 2
13800 företagsfusioner 1
13801 företagsförvärv 1
13802 företagsgrupper 2
13803 företagsgrupperna 2
13804 företagsinterna 1
13805 företagsjuristernas 2
13806 företagskoncentration 1
13807 företagskonsulter 1
13808 företagsledningen 1
13809 företagsledningens 2
13810 företagslikvidation 1
13811 företagslivet 1
13812 företagsnamn 1
13813 företagsnedläggning 1
13814 företagsnedläggningar 1
13815 företagspolitiken 1
13816 företagsråd 2
13817 företagsrådet 6
13818 företagsrådsdirektivet 1
13819 företagsskapande 1
13820 företagsstadgar 1
13821 företagsstruktur 1
13822 företagsstrukturen 2
13823 företagsstöd 2
13824 företagsstöden 1
13825 företagstalangen 1
13826 företagsutveckling 1
13827 företeelse 1
13828 företeelser 2
13829 företräda 7
13830 företrädandet 1
13831 företrädare 116
13832 företrädaren 4
13833 företrädares 3
13834 företrädarna 17
13835 företrädas 4
13836 företrädd 2
13837 företrädda 6
13838 företrädde 1
13839 företräde 5
13840 företräder 22
13841 företrädesvis 2
13842 företräds 3
13843 företrätt 1
13844 förevisas 1
13845 förevändning 7
13846 förevändningar 1
13847 förevändningen 2
13848 förfader 1
13849 förfall 3
13850 förfalla 1
13851 förfallit 1
13852 förfallna 2
13853 förfalskare 1
13854 förfalskas 5
13855 förfalskning 13
13856 förfalskningar 11
13857 förfalskningsutrustning 1
13858 förfarande 48
13859 förfarandefrågor 1
13860 förfaranden 32
13861 förfarandena 14
13862 förfarandet 46
13863 förfaringssätt 1
13864 förfasade 1
13865 förfasar 1
13866 författa 1
13867 författare 8
13868 författaren 4
13869 författares 1
13870 författarna 1
13871 författarnamnet 1
13872 författarnas 1
13873 författat 4
13874 författats 1
13875 författningar 1
13876 författningen 1
13877 författningsenliga 1
13878 författningsfrågor 1
13879 författningsrätt 1
13880 förfela 1
13881 förfiningsarbete 1
13882 förfjol 1
13883 förflutet 1
13884 förflutna 21
13885 förflutnas 1
13886 förflytta 5
13887 förflyttade 2
13888 förflyttar 2
13889 förflyttats 1
13890 förflyttning 6
13891 förflyttningar 1
13892 förflyttningen 1
13893 förfoga 8
13894 förfogande 31
13895 förfoganderätt 1
13896 förfogar 21
13897 förfront 2
13898 förfrysningsskador 1
13899 förfrågan 5
13900 förfrågningar 3
13901 förfäders 1
13902 förfäktar 1
13903 förfärande 5
13904 förfärlig 1
13905 förfärliga 3
13906 förfärligaste 1
13907 förfärligt 5
13908 förfång 3
13909 förfölja 2
13910 förföljare 1
13911 förföljda 1
13912 förföljde 2
13913 förföljelser 3
13914 förföljelserna 3
13915 förföljer 1
13916 förföljs 3
13917 förförisk 2
13918 förförnyelse 1
13919 förfört 1
13920 förgiftar 1
13921 förgiftning 2
13922 förgiftningen 1
13923 förglömma 2
13924 förglömmas 1
13925 förgrening 1
13926 förgrovande 1
13927 förgrunden 5
13928 förgät-mig-ej-blått 1
13929 förgäves 2
13930 förgångna 2
13931 förgångnas 1
13932 förhalande 1
13933 förhand 8
13934 förhandla 26
13935 förhandlade 1
13936 förhandlande 1
13937 förhandlar 3
13938 förhandlarna 2
13939 förhandlas 3
13940 förhandlat 2
13941 förhandlats 2
13942 förhandling 14
13943 förhandlingar 38
13944 förhandlingarna 54
13945 förhandlingarnas 1
13946 förhandlingen 15
13947 förhandlings- 2
13948 förhandlingsbordet 1
13949 förhandlingsflexibilitet 1
13950 förhandlingsforum 1
13951 förhandlingsförfarande 1
13952 förhandlingsgruppen 1
13953 förhandlingsklimatet 1
13954 förhandlingsmandatet 1
13955 förhandlingsparterna 1
13956 förhandlingspartnerna 1
13957 förhandlingsperiod 1
13958 förhandlingsposition 1
13959 förhandlingsprocess 2
13960 förhandlingsprocessen 3
13961 förhandlingsrunda 1
13962 förhandlingsrundan 3
13963 förhandlingsrundorna 1
13964 förhandlingssammanträde 1
13965 förhandlingssammanträdena 1
13966 förhandlingssammanträdet 1
13967 förhandlingssituation 1
13968 förhandlingsskicklighet 1
13969 förhandlingsärenden 1
13970 förhands- 1
13971 förhandsanmälningar 1
13972 förhandsavgörande 2
13973 förhandsavgöranden 1
13974 förhandsbekräftelse 1
13975 förhandsinformation 1
13976 förhandskontroll 2
13977 förhandskontrollen 2
13978 förhastade 3
13979 förhastar 1
13980 förhastat 2
13981 förhindra 73
13982 förhindrade 1
13983 förhindrande 1
13984 förhindrandet 1
13985 förhindrar 9
13986 förhindras 9
13987 förhindrat 2
13988 förhindrats 1
13989 förhistorisk 1
13990 förhoppning 8
13991 förhoppningar 18
13992 förhoppningen 8
13993 förhoppningsvis 8
13994 förhärligade 1
13995 förhärskande 2
13996 förhålla 1
13997 förhållande 56
13998 förhållanden 46
13999 förhållandena 14
14000 förhållandet 30
14001 förhållandevis 3
14002 förhåller 7
14003 förhållit 1
14004 förhållningssätt 4
14005 förhållningssättet 2
14006 förhånas 1
14007 förhöjt 1
14008 förhöll 1
14009 förhörd 1
14010 förintas 1
14011 förintelse 1
14012 förintelsekonferensen 1
14013 förintelsen 2
14014 förirra 1
14015 förkasta 5
14016 förkastade 7
14017 förkastades 3
14018 förkastandet 1
14019 förkastar 9
14020 förkastas 3
14021 förkastat 1
14022 förkastats 2
14023 förkastligt 2
14024 förklara 36
14025 förklarade 24
14026 förklarar 96
14027 förklaras 9
14028 förklarat 12
14029 förklarats 5
14030 förklaring 19
14031 förklaringar 6
14032 förklaringarna 5
14033 förklaringen 4
14034 förklarliga 1
14035 förkläde 1
14036 förkläden 1
14037 förklädet 1
14038 förklädnad 1
14039 förknippad 2
14040 förknippade 5
14041 förknippas 1
14042 förkorta 3
14043 förkortad 1
14044 förkortade 3
14045 förkortas 2
14046 förkortat 1
14047 förkortning 1
14048 förkortningen 1
14049 förkovran 1
14050 förkromade 1
14051 förkrossande 1
14052 förkunna 1
14053 förkunnade 1
14054 förkunnar 1
14055 förkunnat 1
14056 förkunnats 1
14057 förkämpe 3
14058 förkänsla 1
14059 förlagen 1
14060 förlagor 2
14061 förledas 1
14062 förlegad 1
14063 förlegade 1
14064 förlika 1
14065 förlikar 1
14066 förlikning 13
14067 förlikningar 1
14068 förlikningen 13
14069 förliknings- 1
14070 förlikningsetappen 1
14071 förlikningsförfarande 5
14072 förlikningsförfarandet 9
14073 förlikningskommitté 1
14074 förlikningskommittén 11
14075 förlikningskommitténs 6
14076 förlikningsprocess 3
14077 förlikningsprocessen 2
14078 förlikningsvävnad 1
14079 förlisning 7
14080 förlisningen 3
14081 förliste 2
14082 förlita 8
14083 förlitar 8
14084 förloppet 1
14085 förlora 19
14086 förlorad 4
14087 förlorade 13
14088 förlorades 1
14089 förlorar 15
14090 förlorare 1
14091 förloras 1
14092 förlorat 30
14093 förlorats 1
14094 förlossningskliniker 1
14095 förlust 8
14096 förlustbringande 1
14097 förlusten 6
14098 förluster 13
14099 förlusterna 3
14100 förlutet 1
14101 förlägenhet 1
14102 förläggas 1
14103 förläggning 2
14104 förlänga 7
14105 förlängas 2
14106 förlängde 1
14107 förlänger 2
14108 förlängning 9
14109 förlängningen 4
14110 förlängs 4
14111 förlängts 2
14112 förlåt 1
14113 förlåta 2
14114 förlåten 1
14115 förlåter 1
14116 förlöjligar 1
14117 förlöper 1
14118 förmanad 1
14119 förmaning 1
14120 förmedla 9
14121 förmedlade 1
14122 förmedlande 1
14123 förmedlar 2
14124 förmedlare 1
14125 förmedlas 1
14126 förmedling 1
14127 förmenande 3
14128 förment 1
14129 förmenta 2
14130 förmiddag 8
14131 förmiddagen 3
14132 förmiddagens 2
14133 förmiddags 9
14134 förmildrande 1
14135 förmodade 2
14136 förmodar 7
14137 förmodas 1
14138 förmodligen 39
14139 förmyndarskap 1
14140 förmå 9
14141 förmåga 43
14142 förmågan 5
14143 förmån 44
14144 förmånen 1
14145 förmåner 7
14146 förmånligt 1
14147 förmånsavtalen 1
14148 förmånsbehandling 2
14149 förmånspaketet 1
14150 förmånstagare 1
14151 förmånstagarna 1
14152 förmånstillträde 1
14153 förmånsursprung 1
14154 förmår 2
14155 förmås 1
14156 förmått 3
14157 förmögen 1
14158 förmögna 1
14159 förmörkelsen 1
14160 förnamn 1
14161 förnedrande 2
14162 förnedring 1
14163 förneka 11
14164 förnekande 1
14165 förnekar 3
14166 förnekas 4
14167 förnekat 1
14168 förnuft 4
14169 förnuftet 4
14170 förnuftig 10
14171 förnuftiga 10
14172 förnuftigare 2
14173 förnuftigt 16
14174 förnufts- 1
14175 förnumstigt 1
14176 förnya 11
14177 förnyad 1
14178 förnyade 5
14179 förnyande 1
14180 förnyandet 1
14181 förnyar 1
14182 förnyas 2
14183 förnyat 1
14184 förnybar 8
14185 förnybara 40
14186 förnyelse 18
14187 förnyelsen 6
14188 förnyelseområden 1
14189 förnämlig 1
14190 förnämsta 2
14191 förnärma 1
14192 förnärmade 1
14193 förolämpade 1
14194 förolämpande 3
14195 förolämpar 2
14196 förolämpas 1
14197 förolämpat 1
14198 förolämpning 3
14199 förorda 1
14200 förordar 5
14201 förordas 1
14202 förordna 1
14203 förordnanden 1
14204 förordnas 1
14205 förordning 88
14206 förordningar 16
14207 förordningarna 3
14208 förordningen 46
14209 förordningens 6
14210 förorena 2
14211 förorenad 1
14212 förorenade 3
14213 förorenande 10
14214 förorenar 19
14215 förorenare 2
14216 förorenaren 22
14217 förorenarens 3
14218 förorenarna 1
14219 förorenarnas 1
14220 förorenas 5
14221 förorenat 4
14222 förorenats 1
14223 förorening 15
14224 föroreningar 26
14225 föroreningarna 6
14226 föroreningarnas 1
14227 föroreningen 6
14228 föroreningsminskningar 1
14229 förorsaka 3
14230 förorsakad 1
14231 förorsakade 2
14232 förorsakar 2
14233 förorsakas 1
14234 förorsakat 3
14235 förorsakats 3
14236 förorter 5
14237 förorters 1
14238 förpackat 1
14239 förpackning 3
14240 förpackningar 1
14241 förpackningsdirektivet 1
14242 förpassa 2
14243 förpassade 1
14244 förpassades 1
14245 förpassas 1
14246 förpestade 1
14247 förpliktad 1
14248 förpliktade 3
14249 förpliktande 1
14250 förpliktar 3
14251 förpliktas 1
14252 förpliktelse 6
14253 förpliktelsen 3
14254 förpliktelser 14
14255 förpliktiga 1
14256 förpliktigad 2
14257 förpliktigade 2
14258 förpliktigande 1
14259 förpliktigar 1
14260 förpliktigas 1
14261 förpliktigat 3
14262 förr 15
14263 förra 119
14264 förre 6
14265 förresten 5
14266 förrgår 5
14267 förringa 2
14268 förringar 1
14269 förräderi 2
14270 förrädisk 1
14271 förrän 24
14272 förrättar 1
14273 förrättas 1
14274 förråd 1
14275 förrådde 1
14276 förs 18
14277 församlade 1
14278 församling 25
14279 församlingar 3
14280 församlingarna 2
14281 församlingen 27
14282 församlingens 2
14283 församlings 1
14284 försatt 2
14285 förse 18
14286 förseglad 2
14287 försena 4
14288 försenad 8
14289 försenade 7
14290 försenades 1
14291 försenar 1
14292 försenas 2
14293 försenat 5
14294 försening 7
14295 förseningar 8
14296 förseningarna 1
14297 förseningen 6
14298 förser 3
14299 förses 5
14300 försett 2
14301 försetts 1
14302 försiggick 1
14303 försiktig 7
14304 försiktiga 17
14305 försiktighet 14
14306 försiktigheten 2
14307 försiktighetsprincipen 58
14308 försiktighetsprinipen 1
14309 försiktighetsåtgärd 2
14310 försiktighetsåtgärden 1
14311 försiktighetsåtgärder 3
14312 försiktigt 7
14313 försjunken 1
14314 försjunket 1
14315 försjönk 1
14316 förskansad 1
14317 förskingra 1
14318 förskingrat 1
14319 förskingring 2
14320 förskjutas 1
14321 förskjutning 3
14322 förskolor 1
14323 förskonade 1
14324 förskottsbetalningar 1
14325 förskräcka 1
14326 förskräckande 1
14327 förskräcklig 2
14328 förskräckliga 1
14329 förskräckligt 1
14330 förskräckt 2
14331 förskräckta 1
14332 förslag 587
14333 förslagen 42
14334 förslaget 188
14335 förslagets 2
14336 förslagits 2
14337 förslagna 2
14338 förslagsdel 1
14339 förslagspaket 1
14340 förslagsstadiet 1
14341 förslagsställandet 1
14342 förslagsställaren 1
14343 förslavade 1
14344 förslår 2
14345 förslås 2
14346 förslösat 1
14347 försona 3
14348 försonande 3
14349 försoning 8
14350 försoningen 2
14351 försoningshandling 1
14352 försoningskommission 1
14353 försoningsprocessen 1
14354 försoningsprogrammet 2
14355 försonlig 1
14356 förspilla 1
14357 försprång 1
14358 först 144
14359 första 594
14360 förstabehandling 1
14361 förstabehandlingen 2
14362 förstainstansrätt 2
14363 förstainstansrätten 16
14364 förstainstansrättens 3
14365 förstaklasspelare 1
14366 förste 4
14367 förstesekreteraren 1
14368 förstfödde 1
14369 förstklassig 1
14370 förstklassigt 1
14371 förstnämndas 1
14372 förstod 15
14373 förströdd 1
14374 förstulet 1
14375 förställer 1
14376 förställningskonsten 1
14377 förstärka 31
14378 förstärkande 1
14379 förstärkas 7
14380 förstärker 2
14381 förstärkning 15
14382 förstärks 7
14383 förstärkt 11
14384 förstärkta 3
14385 förstå 60
14386 förståeliga 1
14387 förståeligt 5
14388 förståelse 27
14389 förståelsen 2
14390 förstånd 1
14391 förståndiga 2
14392 förstår 75
14393 förstås 21
14394 förstått 22
14395 förstör 18
14396 förstöra 7
14397 förstöras 3
14398 förstörd 1
14399 förstörda 3
14400 förstörde 1
14401 förstördes 4
14402 förstörelse 5
14403 förstörelsen 7
14404 förstöringen 1
14405 förstörs 7
14406 förstört 4
14407 förstörts 9
14408 försumbar 1
14409 försumlighet 1
14410 försumma 1
14411 försummade 1
14412 försummar 2
14413 försummas 1
14414 försummat 1
14415 försummelse 4
14416 försummelsen 1
14417 försummelser 2
14418 försvaga 8
14419 försvagad 1
14420 försvagade 3
14421 försvagades 1
14422 försvagar 7
14423 försvagas 8
14424 försvagats 2
14425 försvagning 3
14426 försvann 12
14427 försvar 31
14428 försvara 43
14429 försvarade 4
14430 försvarades 1
14431 försvarar 18
14432 försvarare 7
14433 försvaras 6
14434 försvarat 10
14435 försvarbara 2
14436 försvaret 11
14437 försvarets 1
14438 försvars- 2
14439 försvarsadvokat 1
14440 försvarsanslag 1
14441 försvarsbeslut 1
14442 försvarsbesparingar 1
14443 försvarsbudgetarna 1
14444 försvarsbudgeten 1
14445 försvarsfrågor 2
14446 försvarshållningen 1
14447 försvarsidentitet 2
14448 försvarsidentiteten 2
14449 försvarsindustrin 1
14450 försvarsinstinkt 1
14451 försvarskapacitet 1
14452 försvarskapaciteten 1
14453 försvarskostnader 1
14454 försvarslösa 2
14455 försvarsmaktens 1
14456 försvarsmedel 1
14457 försvarsminister 2
14458 försvarsministermöte 1
14459 försvarsministern 3
14460 försvarsministrarna 2
14461 försvarsministrarnas 1
14462 försvarsområdet 1
14463 försvarspolitik 18
14464 försvarspolitiken 6
14465 försvarsstrukturer 1
14466 försvarsstyrkor 1
14467 försvarsuppgifter 1
14468 försvarsuppgifterna 1
14469 försvarsutgifter 2
14470 försvarsutvecklingsarbete 1
14471 försvinna 11
14472 försvinnande 4
14473 försvinner 30
14474 försvunnen 1
14475 försvunnit 9
14476 försvåra 2
14477 försvårande 1
14478 försvårar 3
14479 försvåras 3
14480 försäkra 41
14481 försäkrade 7
14482 försäkran 2
14483 försäkrar 7
14484 försäkrats 1
14485 försäkring 1
14486 försäkringar 9
14487 försäkringarna 1
14488 försäkringsavgifter 1
14489 försäkringsbedrägerier 1
14490 försäkringsbevis 3
14491 försäkringsbolag 2
14492 försäkringsbolagen 1
14493 försäkringsbolaget 1
14494 försäkringsmarknaden 1
14495 försäkringsrättigheter 1
14496 försäkringssektorn 1
14497 försäkringsskydd 2
14498 försäkringssystem 1
14499 försäkringssystemen 1
14500 försäljare 1
14501 försäljaren 2
14502 försäljning 9
14503 försäljningen 2
14504 försäljningsnedgången 2
14505 försäljningsrapport 1
14506 försäljningsrapporten 1
14507 försäljningsvolym 1
14508 försäljs 1
14509 försämra 5
14510 försämrad 3
14511 försämrade 4
14512 försämrande 1
14513 försämras 6
14514 försämring 4
14515 försämringar 1
14516 försämringarna 1
14517 försämringen 3
14518 försändelserna 1
14519 försänkts 1
14520 försätter 1
14521 försåg 2
14522 försågs 1
14523 försåtligt 1
14524 försåvitt 1
14525 försök 32
14526 försöka 108
14527 försöken 4
14528 försöker 78
14529 försöket 3
14530 försökslaboratorium 1
14531 försöksmässigt 1
14532 försökt 24
14533 försökte 43
14534 försökts 1
14535 försörja 3
14536 försörjer 1
14537 försörjning 4
14538 försörjningsgrund 1
14539 fört 13
14540 förtal 1
14541 förtecken 1
14542 förtecknades 1
14543 förteckning 7
14544 förteckningen 8
14545 förtennad 1
14546 förtid 1
14547 förtida 1
14548 förtidspension 2
14549 förtidspensionerade 2
14550 förtidspensionering 2
14551 förtidspensioneringssystemet 2
14552 förtjusande 1
14553 förtjusning 3
14554 förtjust 4
14555 förtjusta 2
14556 förtjäna 4
14557 förtjänade 2
14558 förtjänar 41
14559 förtjänats 1
14560 förtjänst 2
14561 förtjänsten 2
14562 förtjänster 3
14563 förtjänstfulla 1
14564 förtjänstfullt 2
14565 förtjänt 1
14566 förtjänta 2
14567 förtroende 67
14568 förtroendeförskott 1
14569 förtroendeklyftan 1
14570 förtroendekris 2
14571 förtroenden 1
14572 förtroendeposter 1
14573 förtroenderöst 1
14574 förtroendeskapande 3
14575 förtroendet 17
14576 förtroendeuppbyggnaden 1
14577 förtroendevald 4
14578 förtroendevalda 2
14579 förtroendeväckande 1
14580 förtrogen 1
14581 förtrogna 1
14582 förtrollar 1
14583 förtrollat 1
14584 förtryck 4
14585 förtryckande 2
14586 förtryckare 1
14587 förtryckarhierarki 1
14588 förtryckarregimen 1
14589 förtrycket 2
14590 förtrycktas 1
14591 förtrytelse 1
14592 förträffliga 2
14593 förträfflighet 1
14594 förtränger 1
14595 förts 12
14596 förtursbehandling 1
14597 förtvivla 1
14598 förtvivlade 3
14599 förtvivlan 6
14600 förtvivlat 2
14601 förtydliga 6
14602 förtydligande 2
14603 förtydliganden 4
14604 förtäckt 2
14605 förtäckta 2
14606 förtära 1
14607 förtärande 1
14608 förtätad 1
14609 förtöjd 1
14610 förtöjda 1
14611 förunderligt 2
14612 förundersökningshandlingar 1
14613 förundra 1
14614 förundran 1
14615 förut 12
14616 förutan 1
14617 förutbestämd 1
14618 förutbestämt 1
14619 förutom 44
14620 förutsatt 3
14621 förutsatte 1
14622 förutse 6
14623 förutsebar 1
14624 förutsedd 1
14625 förutseende 2
14626 förutser 1
14627 förutses 5
14628 förutsett 2
14629 förutsetts 3
14630 förutspå 1
14631 förutspåddes 2
14632 förutspås 1
14633 förutsäga 3
14634 förutsägbar 2
14635 förutsägbara 1
14636 förutsägbart 1
14637 förutsägelse 2
14638 förutsätta 2
14639 förutsättas 1
14640 förutsätter 30
14641 förutsättning 39
14642 förutsättningar 24
14643 förutsättningarna 11
14644 förutsättningen 4
14645 förutsättningslös 1
14646 förutsätts 1
14647 förutvarande 3
14648 förvalta 11
14649 förvaltad 2
14650 förvaltande 1
14651 förvaltar 4
14652 förvaltare 2
14653 förvaltaren 2
14654 förvaltas 4
14655 förvaltning 62
14656 förvaltningar 6
14657 förvaltningarna 2
14658 förvaltningarnas 1
14659 förvaltningen 36
14660 förvaltningens 1
14661 förvaltningsbolag 6
14662 förvaltningsbolagen 3
14663 förvaltningsbolaget 1
14664 förvaltningsförfarande 3
14665 förvaltningsförfaranden 1
14666 förvaltningsförfarandet 3
14667 förvaltningskommittéer 1
14668 förvaltningskostnaderna 2
14669 förvaltningsmyndigheters 1
14670 förvaltningsområde 1
14671 förvaltningsorgan 1
14672 förvaltningsprinciper 1
14673 förvaltningsrätt 2
14674 förvaltningssed 1
14675 förvaltningsstrukturen 1
14676 förvaltningssystem 3
14677 förvaltningstekniska 1
14678 förvaltningsuppdrag 1
14679 förvaltningsuppgifterna 1
14680 förvaltningsverksamhet 1
14681 förvaltningsåtgärder 1
14682 förvaltningsåtgärderna 1
14683 förvandla 6
14684 förvandlade 1
14685 förvandlar 5
14686 förvandlas 8
14687 förvandlat 1
14688 förvandlats 4
14689 förvanskar 1
14690 förvanskas 1
14691 förvanskats 1
14692 förvar 1
14693 förvaras 1
14694 förvarna 1
14695 förvarnade 1
14696 förvarningssystem 1
14697 förverkliga 23
14698 förverkligades 1
14699 förverkligande 1
14700 förverkligandet 6
14701 förverkligas 13
14702 förverkligats 4
14703 förvirrad 3
14704 förvirrade 2
14705 förvirrande 2
14706 förvirrar 1
14707 förvirrat 2
14708 förvirring 13
14709 förvirringen 1
14710 förvisade 1
14711 förvisats 2
14712 förvisningsorder 1
14713 förvissad 2
14714 förvissade 1
14715 förvissning 1
14716 förvisso 24
14717 förvriden 2
14718 förvränga 1
14719 förvrängd 1
14720 förväg 21
14721 förvägra 2
14722 förvägrad 1
14723 förvägrades 2
14724 förvägrar 2
14725 förvägras 1
14726 förvägrats 2
14727 förvänta 10
14728 förväntade 2
14729 förväntades 2
14730 förväntan 2
14731 förväntar 45
14732 förväntas 7
14733 förväntat 6
14734 förväntningar 20
14735 förväntningarna 5
14736 förvärra 2
14737 förvärrade 1
14738 förvärras 5
14739 förvärrat 2
14740 förvärrats 3
14741 förvärva 4
14742 förvärvas 1
14743 förvärvat 1
14744 förvärvsarbete 4
14745 förvärvsarbetet 2
14746 förväxla 2
14747 förväxlar 1
14748 förvåna 2
14749 förvånad 7
14750 förvånade 3
14751 förvånande 3
14752 förvånansvärt 3
14753 förvånar 2
14754 förvånas 2
14755 förvånats 1
14756 förvåning 5
14757 förädla 2
14758 förädlade 2
14759 förälder 1
14760 föräldraledighet 2
14761 föräldrar 15
14762 föräldrarnas 1
14763 föräldrars 3
14764 förälskad 1
14765 föränderliga 3
14766 förändra 27
14767 förändrade 4
14768 förändrades 5
14769 förändrar 6
14770 förändras 22
14771 förändrat 3
14772 förändrats 8
14773 förändring 42
14774 förändringar 65
14775 förändringarna 14
14776 förändringen 3
14777 förändringens 1
14778 förändringsarbetet 2
14779 förändringsprocesser 1
14780 föråldrad 1
14781 föråldrade 10
14782 föråldrat 2
14783 förödande 11
14784 förödelse 3
14785 förödmjukande 1
14786 förödmjukelser 1
14787 förökar 1
14788 förökning 1
14789 förövades 1
14790 förövaren 2
14791 förövarna 2
14792 föröver 1
14793 fötter 12
14794 fötterna 7
14795 fötts 2
14796 g 3
14797 gaberdin 1
14798 gaffel 3
14799 gaffeldukar 1
14800 gaffeln 1
14801 gafflarnas 1
14802 gagn 4
14803 gagna 1
14804 gagnar 3
14805 gagnat 2
14806 galakvinnor 1
14807 galax 1
14808 galaxer 1
14809 galen 5
14810 galenskap 1
14811 galenskapen 1
14812 galenskaps 1
14813 galiciska 1
14814 galjonsfiguren 1
14815 galleon 1
14816 galler 2
14817 gallerstängerna 2
14818 gallren 1
14819 gallret 2
14820 gallring 1
14821 gallringen 1
14822 galna 5
14823 galning 1
14824 galningar 2
14825 galopp 1
14826 galopperande 1
14827 gamla 99
14828 gamle 5
14829 gammal 28
14830 gammaldags 1
14831 gammalmodig 1
14832 gammalt 8
14833 gangstertyper 1
14834 ganska 96
14835 gapade 1
14836 gapet 1
14837 gapskratt 2
14838 garage 1
14839 garant 6
14840 garantera 116
14841 garanterad 2
14842 garanterade 4
14843 garanterar 31
14844 garanteras 13
14845 garanterat 6
14846 garanterats 1
14847 garanti 20
14848 garantier 30
14849 garantierna 9
14850 garantifonden 3
14851 garantin 5
14852 garantisektion 1
14853 garantisektionen 1
14854 garantisystemet 1
14855 garde-länderna 2
14856 garderobsdörren 1
14857 gardinen 1
14858 garn 1
14859 gas 2
14860 gaskammare 1
14861 gassade 1
14862 gasutsläpp 1
14863 gata 3
14864 gatan 25
14865 gathörn 1
14866 gathörnstyper 1
14867 gator 4
14868 gatorna 6
14869 gatornas 1
14870 gav 79
14871 gavel 2
14872 gavs 10
14873 gazatska 1
14874 ge 411
14875 gedigen 1
14876 gediget 1
14877 gedigna 2
14878 gehör 2
14879 gelikar 1
14880 gemener 3
14881 gemensam 140
14882 gemensamma 391
14883 gemensamt 57
14884 gemenskap 23
14885 gemenskapen 129
14886 gemenskapens 184
14887 gemenskaper 1
14888 gemenskaperna 5
14889 gemenskapernas 8
14890 gemenskaplig 1
14891 gemenskaps- 1
14892 gemenskapsarvet 1
14893 gemenskapsaspekt 1
14894 gemenskapsavtal 1
14895 gemenskapsbefogenheterna 1
14896 gemenskapsbestämmelser 2
14897 gemenskapsbestämmelserna 3
14898 gemenskapsbidrag 1
14899 gemenskapsbidraget 1
14900 gemenskapsbudgeten 5
14901 gemenskapsdimensionen 1
14902 gemenskapsdirektiv 2
14903 gemenskapsdirektiven 2
14904 gemenskapsengagemang 1
14905 gemenskapsfilosofin 1
14906 gemenskapsfond 2
14907 gemenskapsfonder 1
14908 gemenskapsfrågor 1
14909 gemenskapsfördragens 1
14910 gemenskapsgrupper 2
14911 gemenskapshamnar 1
14912 gemenskapshamnarna 1
14913 gemenskapshamnarnas 1
14914 gemenskapsinförlivande 1
14915 gemenskapsinitiativ 20
14916 gemenskapsinitiativen 13
14917 gemenskapsinitiativet 26
14918 gemenskapsinitiativets 1
14919 gemenskapsinitiativs 1
14920 gemenskapsinsatserna 1
14921 gemenskapsinstitutionerna 4
14922 gemenskapsinstitutionernas 3
14923 gemenskapsinstrument 3
14924 gemenskapsintresse 1
14925 gemenskapsintressen 1
14926 gemenskapskonstruktion 1
14927 gemenskapskontroll 1
14928 gemenskapslag 1
14929 gemenskapslagstiftning 5
14930 gemenskapslagstiftningen 13
14931 gemenskapslagstiftningens 1
14932 gemenskapsmaskinen 1
14933 gemenskapsmaskinens 1
14934 gemenskapsmedborgare 1
14935 gemenskapsnivå 28
14936 gemenskapsnormerna 1
14937 gemenskapsområdet 1
14938 gemenskapsorgan 2
14939 gemenskapspelaren 3
14940 gemenskapsplanet 1
14941 gemenskapspolitik 5
14942 gemenskapspolitiken 6
14943 gemenskapspolitikens 2
14944 gemenskapspreferensen 1
14945 gemenskapsprocessen 1
14946 gemenskapsproduktionen 1
14947 gemenskapsprogram 5
14948 gemenskapsprogrammen 5
14949 gemenskapsprogrammet 1
14950 gemenskapsram 2
14951 gemenskapsramen 1
14952 gemenskapsregister 1
14953 gemenskapsregler 2
14954 gemenskapsreglerna 5
14955 gemenskapsresurserna 2
14956 gemenskapsrätt 1
14957 gemenskapsrätten 17
14958 gemenskapsstadga 1
14959 gemenskapsstrategi 1
14960 gemenskapsstrukturerna 1
14961 gemenskapsstöd 2
14962 gemenskapsstödets 1
14963 gemenskapsstödramar 1
14964 gemenskapsstödramarna 1
14965 gemenskapsstödramen 11
14966 gemenskapssystem 1
14967 gemenskapstexter 1
14968 gemenskapsvatten 2
14969 gemenskapsvattnen 1
14970 gemenskapsåtgärd 1
14971 gemenskapsåtgärder 6
14972 gement 1
14973 gemyt 1
14974 gemål 1
14975 genant 1
14976 genast 24
14977 gender 7
14978 genderkurser 1
14979 genderutbildning 1
14980 genderutbildningen 1
14981 genera 1
14982 generad 3
14983 generade 1
14984 general 4
14985 generaladvokaten 1
14986 generalangrepp 1
14987 generaldirektorat 10
14988 generaldirektoraten 3
14989 generaldirektoratet 9
14990 generaldirektör 2
14991 generaldirektören 1
14992 generaldirektörens 1
14993 generaler 1
14994 generalförsamling 1
14995 generalförsamlingen 2
14996 generalisera 1
14997 generaliserade 1
14998 generaliseras 1
14999 generaliseringar 1
15000 generalklausul 1
15001 generalsekretariat 1
15002 generalsekreterare 22
15003 generalsekreteraren 3
15004 generalsekreterares 2
15005 generande 2
15006 generation 2
15007 generationen 2
15008 generationer 11
15009 generationerna 2
15010 generationernas 2
15011 generationers 1
15012 generell 8
15013 generella 9
15014 generellt 12
15015 generera 4
15016 genererar 7
15017 genereras 1
15018 generiska 1
15019 generositet 3
15020 generositeten 1
15021 generös 4
15022 generösa 2
15023 generösare 1
15024 generöst 3
15025 genetiskt 25
15026 gengäld 5
15027 gengångare 1
15028 geni 1
15029 genial 1
15030 genier 1
15031 genljud 1
15032 genmodifieringsteknik 1
15033 genom 708
15034 genomarbetad 1
15035 genomarbetat 2
15036 genomblickbar 2
15037 genomblickbarhet 5
15038 genomblickbarheten 1
15039 genomblickbart 3
15040 genomblåstes 1
15041 genombrott 5
15042 genombrottet 1
15043 genomdriva 6
15044 genomdrivande 1
15045 genomdrivit 1
15046 genomdrivs 2
15047 genomfarter 1
15048 genomför 18
15049 genomföra 144
15050 genomförande 34
15051 genomförandebefogenheter 4
15052 genomförandebeslut 1
15053 genomförandebestämmelserna 1
15054 genomförandeförordningarna 1
15055 genomföranden 1
15056 genomförandena 1
15057 genomförandet 76
15058 genomförandeverksamheterna 1
15059 genomförandeåtgärd 1
15060 genomförandeåtgärden 2
15061 genomförandeåtgärder 3
15062 genomföras 55
15063 genomförbar 5
15064 genomförbara 4
15065 genomförbarhet 2
15066 genomförbarheten 1
15067 genomförbart 5
15068 genomförd 4
15069 genomförda 3
15070 genomförde 5
15071 genomfördes 9
15072 genomförs 39
15073 genomfört 8
15074 genomförts 18
15075 genomgick 3
15076 genomgripande 16
15077 genomgå 5
15078 genomgående 3
15079 genomgång 5
15080 genomgången 1
15081 genomgår 5
15082 genomgått 7
15083 genomled 1
15084 genomlidandet 1
15085 genomläsning 3
15086 genomskinliga 2
15087 genomskinligt 1
15088 genomslag 4
15089 genomslagskraft 2
15090 genomsnitt 12
15091 genomsnittet 6
15092 genomsnittlig 4
15093 genomsnittliga 5
15094 genomsnittligen 1
15095 genomsnittligt 1
15096 genomsnittsregionerna 1
15097 genomströmmar 1
15098 genomsynlighet 1
15099 genomsyra 4
15100 genomsyrade 1
15101 genomsyrar 1
15102 genomsyras 2
15103 genomsyrats 1
15104 genomsöks 1
15105 genomsökte 1
15106 genomträngande 2
15107 genomträngning 1
15108 genomtänkt 1
15109 genomtänkta 1
15110 gensvar 2
15111 gentemot 78
15112 gentjänster 1
15113 genuin 2
15114 genusdimensionen 1
15115 geografisk 5
15116 geografiska 20
15117 geografiskt 5
15118 geologiska 1
15119 geologiskt 1
15120 geometri 1
15121 geopolitiska 2
15122 geostrategiska 3
15123 geostrategiskt 1
15124 ger 224
15125 gerillamönstret 1
15126 ges 46
15127 gest 12
15128 gestalt 1
15129 gestalta 1
15130 gester 1
15131 gesterna 1
15132 gestikulerade 1
15133 gestikulerande 1
15134 geting 1
15135 gett 69
15136 getter 2
15137 getton 2
15138 getts 2
15139 gevär 1
15140 geväret 1
15141 ghananer 1
15142 ghetto 1
15143 ghoulen 1
15144 gick 132
15145 gift 3
15146 gifta 2
15147 giftblandningarna 1
15148 gifte 4
15149 giftig 1
15150 giftiga 6
15151 giftigt 1
15152 giftkatastrof 1
15153 giftutsläppet 1
15154 gigantisk 3
15155 gigantiska 4
15156 gigantiskt 1
15157 giljotinen 1
15158 gilla 4
15159 gillade 4
15160 gillades 1
15161 gillande 3
15162 gillar 6
15163 gillat 1
15164 gillrat 1
15165 giltig 5
15166 giltiga 2
15167 giltighet 6
15168 giltigheten 3
15169 giltighetstid 11
15170 giltighetstiden 3
15171 giltigt 3
15172 gin 4
15173 ginge 1
15174 giromedel 1
15175 gissa 5
15176 gissade 2
15177 gisslan 5
15178 gitarrer 1
15179 givande 3
15180 givandet 1
15181 givare 9
15182 givares 1
15183 givarkonferensen 1
15184 givarlandens 1
15185 givarlandet 1
15186 givarländer 1
15187 givarländerna 2
15188 givarna 6
15189 givarnas 1
15190 givarsamfundet 1
15191 givas 1
15192 given 2
15193 gives 1
15194 givet 3
15195 givetvis 72
15196 givit 12
15197 givits 2
15198 givmild 1
15199 givna 3
15200 gjord 3
15201 gjorda 1
15202 gjorde 119
15203 gjordes 17
15204 gjort 208
15205 gjorts 56
15206 glad 56
15207 glada 9
15208 gladde 2
15209 gladeligen 1
15210 glamorös 1
15211 glans 2
15212 glansdager 1
15213 glas 11
15214 glasdörr 1
15215 glasen 1
15216 glaset 1
15217 glashus 1
15218 glasklart 1
15219 glasmonter 1
15220 glasmontrarna 1
15221 glaspärlor 1
15222 glass 2
15223 glassförsäljarnas 1
15224 glasskivorna 1
15225 glasögon 4
15226 glasögonbärare 1
15227 glasögonen 5
15228 glatt 4
15229 gled 6
15230 glesa 1
15231 glesbefolkade 3
15232 glesbygden 1
15233 glesbygdsområden 1
15234 glest 3
15235 glida 1
15236 glider 2
15237 glimma 1
15238 glimmade 3
15239 glimmande 1
15240 glimmar 1
15241 glimt 2
15242 glimtar 1
15243 glimten 1
15244 glitterögd 1
15245 glittrande 4
15246 global 17
15247 globala 30
15248 globaliserad 3
15249 globaliserade 4
15250 globaliserande 1
15251 globalisering 12
15252 globaliseringen 32
15253 globaliseringens 3
15254 globaliseringsdiskussionen 1
15255 globaliseringsprocessen 1
15256 globaliteten 1
15257 globalt 13
15258 glodde 2
15259 glorifiering 1
15260 glunkades 1
15261 glupskhet 1
15262 gläder 58
15263 glädja 14
15264 glädjande 16
15265 glädjas 4
15266 glädje 17
15267 glädjen 1
15268 glädjevitt 1
15269 gläds 12
15270 glänsande 3
15271 glänste 1
15272 glänt 1
15273 glöd 2
15274 glödande 1
15275 glödde 1
15276 glödhög 1
15277 glödlampa 1
15278 glödlampor 1
15279 glöm 1
15280 glömd 1
15281 glömde 7
15282 glömma 44
15283 glömmas 1
15284 glömmer 10
15285 glöms 1
15286 glömska 1
15287 glömskan 1
15288 glömt 9
15289 gnista 1
15290 gnistor 2
15291 gnistrade 1
15292 gnistrande 1
15293 gnistregnet 1
15294 gnome 1
15295 gnomehålen 1
15296 gnomen 1
15297 gnomens 1
15298 gnomer 3
15299 gnuggar 1
15300 gnutta 2
15301 gnäller 1
15302 gnället 1
15303 goals 2
15304 god 66
15305 goda 98
15306 godafton 1
15307 godas 1
15308 gode 2
15309 godhet 1
15310 godhjärtad 1
15311 godkänd 5
15312 godkända 8
15313 godkände 20
15314 godkändes 11
15315 godkänna 49
15316 godkännande 30
15317 godkännandeförbehåll 1
15318 godkännandena 1
15319 godkännandet 9
15320 godkännas 18
15321 godkänner 29
15322 godkänns 4
15323 godkänt 21
15324 godkänts 22
15325 godmodigt 1
15326 godo 5
15327 gods 39
15328 godset 1
15329 godsets 1
15330 godsfinka 1
15331 godstransporter 1
15332 godstransporterna 1
15333 godta 24
15334 godtagbar 9
15335 godtagbara 7
15336 godtagbart 17
15337 godtagit 3
15338 godtagits 1
15339 godtar 15
15340 godtas 11
15341 godtog 4
15342 godtogs 3
15343 godtycke 1
15344 godtycklig 2
15345 godtyckliga 2
15346 godtyckligt 4
15347 gojernas 1
15348 golfförsäljningen 2
15349 golliwog 1
15350 golvet 8
15351 gom 1
15352 good 3
15353 gossarna 1
15354 gosse 1
15355 gossen 1
15356 gott 50
15357 gottgöra 2
15358 gottgörelse 1
15359 gottgörelsen 1
15360 governance 5
15361 government 1
15362 governments 1
15363 governo 2
15364 grabb 1
15365 gracila 1
15366 graciös 1
15367 grad 62
15368 graden 5
15369 grader 9
15370 graderna 1
15371 gradvis 16
15372 gradvisa 4
15373 gradvist 1
15374 graecas 1
15375 grafiskt 1
15376 gram 4
15377 grammatikstruktur 1
15378 grammofonnål 1
15379 grammofonskivor 1
15380 granadillpuddingen 1
15381 granaterna 1
15382 grand 6
15383 grannar 12
15384 granne 1
15385 grannförbindelser 1
15386 grannlagenhet 1
15387 grannland 1
15388 grannlandet 2
15389 grannländer 4
15390 grannländerna 9
15391 grannländernas 1
15392 grannregioner 1
15393 grannregionernas 1
15394 grannskap 2
15395 grannskapet 2
15396 grannsämja 1
15397 grannsämjan 1
15398 granska 44
15399 granskade 7
15400 granskades 1
15401 granskar 10
15402 granskas 14
15403 granskat 3
15404 granskats 3
15405 granskning 31
15406 granskningar 1
15407 granskningarna 2
15408 granskningen 9
15409 granskningsenhet 1
15410 granskningsmekanismer 1
15411 granskningsprocess 3
15412 granskningssystemet 1
15413 gras 1
15414 gras-fest 1
15415 gras-fester 1
15416 gratis 12
15417 gratulationer 8
15418 gratulera 64
15419 gratulerade 1
15420 gratulerar 21
15421 gratulerat 1
15422 grav 3
15423 grava 1
15424 gravar 3
15425 gravarna 1
15426 graverande 4
15427 gravgrottor 1
15428 gravida 3
15429 graviditet 1
15430 graviditetsmånad 1
15431 graviterade 1
15432 gravt 1
15433 gravvalv 1
15434 green 1
15435 grej 1
15436 grejor 1
15437 grek 1
15438 grekcypriotiska 2
15439 grekerna 2
15440 grekisk-turkiska 1
15441 grekiska 28
15442 grekiskt 1
15443 gren 2
15444 grenar 3
15445 grenarna 3
15446 grenen 3
15447 grep 4
15448 grepen 1
15449 grepp 5
15450 greppa 1
15451 greppade 2
15452 greps 2
15453 grevskapsrådet 1
15454 grillad 1
15455 grillade 1
15456 grimas 2
15457 grimaserande 1
15458 grimskaft 2
15459 grina 1
15460 grind 1
15461 gripa 6
15462 gripande 1
15463 gripas 1
15464 griper 3
15465 gripit 2
15466 gripna 1
15467 grips 1
15468 grisfet 1
15469 griskött 1
15470 grisköttssektorn 1
15471 grissinistänger 1
15472 grodor 2
15473 grogrund 1
15474 grogrunden 1
15475 grop 2
15476 groteska 1
15477 group 1
15478 grov 1
15479 grova 1
15480 grovt 1
15481 grund 317
15482 grund- 2
15483 grunda 2
15484 grundad 11
15485 grundade 5
15486 grundades 4
15487 grundandet 2
15488 grundar 24
15489 grundarna 2
15490 grundas 13
15491 grundat 14
15492 grundbegrepp 1
15493 grundbulten 1
15494 grunddokument 2
15495 grunden 60
15496 grundens 1
15497 grunder 13
15498 grunderna 3
15499 grundfördrag 1
15500 grundförståelsen 1
15501 grundförtroende 1
15502 grundförutsättning 2
15503 grundförutsättningar 1
15504 grundidén 1
15505 grundingredienserna 1
15506 grundinställning 2
15507 grundkoncept 2
15508 grundkurs 1
15509 grundlagsstridigt 1
15510 grundlig 6
15511 grundliga 4
15512 grundligare 2
15513 grundligt 13
15514 grundläggande 240
15515 grundläggarna 1
15516 grundorsakerna 1
15517 grundpelare 1
15518 grundpelaren 1
15519 grundprincip 2
15520 grundprincipen 2
15521 grundprinciper 1
15522 grundprinciperna 2
15523 grundproblem 1
15524 grundproblemet 1
15525 grundregeln 1
15526 grundsatsen 3
15527 grundsatserna 1
15528 grundskolan 1
15529 grundskolebarn 1
15530 grundskolorna 1
15531 grundsten 2
15532 grundstenar 1
15533 grundstomme 1
15534 grundstommen 2
15535 grundsyn 1
15536 grundtankarna 1
15537 grundtes 1
15538 grundtonen 1
15539 grundtrygghet 1
15540 grundtryggheten 1
15541 grundutbildning 2
15542 grundval 52
15543 grundvalar 3
15544 grundvalen 2
15545 grundvatten 5
15546 grundvattenakviferer 1
15547 grundvattenförekomsternas 1
15548 grundvattenkvalitet 1
15549 grundvattenkvaliteten 1
15550 grundvattenlagren 1
15551 grundvattenreserverna 2
15552 grundvattenstatus 2
15553 grundvattenstatusen 1
15554 grundvattnet 11
15555 grundvillkor 1
15556 grundämnen 1
15557 grupp 225
15558 gruppen 69
15559 gruppens 10
15560 grupper 81
15561 gruppera 9
15562 grupperade 3
15563 grupperas 1
15564 gruppering 1
15565 grupperingar 4
15566 grupperna 42
15567 gruppernas 1
15568 gruppers 5
15569 gruppkollega 1
15570 gruppkolleger 1
15571 gruppnivå 1
15572 gruppnivåer 2
15573 gruppnivån 2
15574 gruppordförande 1
15575 gruppordförandekommittén 1
15576 grupps 16
15577 grupptillhörighet 2
15578 gruppundantaget 1
15579 gruppvis 1
15580 gruva 3
15581 gruvan 1
15582 gruvarbetarfacket 1
15583 gruvbolaget 1
15584 gruvbolagets 1
15585 gruvbrytningen 1
15586 gruvbrytningens 1
15587 gruvbrytningsföretag 1
15588 gruvjobbarpub 1
15589 gruvkoncessionsföretag 1
15590 gruvnäringen 1
15591 gruvor 2
15592 grym 2
15593 grymhet 1
15594 grymt 6
15595 grymta 1
15596 grytor 1
15597 grytorna 1
15598 grädde 1
15599 gräddtårtan 1
15600 gräl 4
15601 grälade 2
15602 grälar 1
15603 grämelse 1
15604 gränd 1
15605 gränden 2
15606 gräns 9
15607 gränsar 4
15608 gränsdragning 1
15609 gränsen 13
15610 gränser 54
15611 gränserna 39
15612 gränsfrågan 3
15613 gränskonflikter 1
15614 gränskontroll 3
15615 gränskontroller 2
15616 gränskontrollerna 1
15617 gränskontrollorganet 1
15618 gränskontrollsystemet 1
15619 gränslandet 1
15620 gränslinjen 1
15621 gränslöst 2
15622 gränsområde 2
15623 gränsområden 2
15624 gränsområdena 4
15625 gränsområdenas 1
15626 gränsprocesserna 1
15627 gränsregioner 2
15628 gränsregionerna 2
15629 gränsregionernas 1
15630 gränssmugglingen 1
15631 gränssnitt 1
15632 gränsstilen 1
15633 gränssäkerhet 1
15634 gränstrakterna 2
15635 gränsvärde 1
15636 gränsvärdena 1
15637 gränsövergripande 1
15638 gränsövergångsnivå 1
15639 gränsöverskridande 54
15640 gräset 8
15641 gräsligas 1
15642 gräslighet 1
15643 gräsligt 1
15644 gräsmatta 1
15645 gräsmattan 3
15646 gräsrotsgrupper 1
15647 gräsrotsnivå 1
15648 grässkjul 1
15649 grät 2
15650 grävde 1
15651 gräver 2
15652 grävt 1
15653 grå 6
15654 grå- 1
15655 grådaskighet 1
15656 grånad 1
15657 gråt 2
15658 gråta 2
15659 grått 3
15660 gråvita 1
15661 gråzon 2
15662 grödor 1
15663 grön 14
15664 gröna 54
15665 grönare 1
15666 grönas 3
15667 grönbok 1
15668 grönböcker 1
15669 grönfodrad 1
15670 grönsaker-snap 1
15671 grönsakerna 1
15672 grönska 2
15673 grönskande 1
15674 grönt 4
15675 gröt 1
15676 grövsta 2
15677 gubbe 1
15678 gubben 4
15679 gud 3
15680 gudabild 1
15681 gudinna 1
15682 gudmor 1
15683 guds 3
15684 gudskelov 1
15685 gul 2
15686 gula 2
15687 gulag 1
15688 gulblekt 1
15689 gulbruna 1
15690 guld 5
15691 guld-metall 1
15692 guldbokstäver 1
15693 gulden 1
15694 guldet 2
15695 guldgruva 1
15696 guldhöna 1
15697 guldringar 1
15698 guldsandal 1
15699 gullade 1
15700 gullegrisar 1
15701 gult 4
15702 gummidocka 1
15703 gummiparagraf 1
15704 gummistämpel 1
15705 gummistövlar 1
15706 gunga 1
15707 gungade 1
15708 gungades 1
15709 gungande 1
15710 gungar 1
15711 guvenörskap 1
15712 guvernör 3
15713 guvernören 2
15714 guvernörens 1
15715 gyllene 7
15716 gym 1
15717 gymnasiet 1
15718 gymnasium 1
15719 gymnastikskor 1
15720 gynna 15
15721 gynnade 6
15722 gynnar 10
15723 gynnas 1
15724 gynnsam 4
15725 gynnsamma 7
15726 gynnsamt 1
15727 gyroskop 1
15728 gyttjemark 1
15729 gyttjig 1
15730 gyttjiga 1
15731 gäck 1
15732 gäldenärens 1
15733 gälla 47
15734 gällande 61
15735 gällde 24
15736 gäller 1028
15737 gällt 5
15738 gäng 4
15739 gängse 1
15740 gärna 123
15741 gärning 3
15742 gärningar 5
15743 gärningsmannen 1
15744 gärningsmän 2
15745 gäspa 1
15746 gäspade 1
15747 gäss 1
15748 gäst 4
15749 gäster 1
15750 gästerna 2
15751 gästfrihet 1
15752 gästhyddan 1
15753 gästrummet 1
15754 gå 252
15755 gång 256
15756 gångarna 3
15757 gången 85
15758 gånger 87
15759 gångna 8
15760 gångs 5
15761 går 318
15762 gård 1
15763 gårdagens 9
15764 gårdar 1
15765 gården 4
15766 gås 2
15767 gåsmarsch 1
15768 gåspenna 1
15769 gåta 4
15770 gåtan 1
15771 gåtfulla 1
15772 gåtfullt 2
15773 gått 67
15774 gåva 1
15775 göda 1
15776 gödsel 1
15777 gödseln 1
15778 gömda 1
15779 gömde 1
15780 gömma 2
15781 gömmas 1
15782 gömmer 5
15783 gömställe 1
15784 gömts 1
15785 gör 399
15786 göra 815
15787 göras 71
15788 görs 50
15789 ha 634
15790 habitat- 1
15791 habitatdirektiv 1
15792 habitatdirektivet 2
15793 hack 1
15794 hackande 1
15795 hade 813
15796 haft 93
15797 hajade 1
15798 haka 1
15799 hakan 1
15800 hakat 1
15801 halka 1
15802 halkade 2
15803 halkar 1
15804 hallen 4
15805 hallickaktigt 1
15806 hallmattan 1
15807 halm 2
15808 halogenerade 1
15809 hals 8
15810 halsar 2
15811 halsarna 1
15812 halsband 1
15813 halsbrytande 1
15814 halsduk 1
15815 halsen 6
15816 halt 2
15817 halta 1
15818 halte 1
15819 halv 12
15820 halva 10
15821 halvan 1
15822 halvdunklet 1
15823 halverades 1
15824 halverats 1
15825 halveringen 1
15826 halvhjärtade 1
15827 halvhjärtat 1
15828 halvideologiska 1
15829 halvkloten 1
15830 halvklädda 1
15831 halvmiljon 1
15832 halvminnen 1
15833 halvoffentliga 1
15834 halvor 1
15835 halvsovit 1
15836 halvt 7
15837 halvtidsbedömningen 1
15838 halvtimme 5
15839 halvvuxen 1
15840 halvvägs 6
15841 halvår 1
15842 halvåret 3
15843 halvårsskifte 1
15844 halvårsskiftet 2
15845 halvö 2
15846 halvön 2
15847 hamburgare 2
15848 hammare 2
15849 hamn 22
15850 hamna 8
15851 hamnade 3
15852 hamnanläggningen 1
15853 hamnar 47
15854 hamnarna 20
15855 hamnarnas 1
15856 hamnat 9
15857 hamnavgiften 2
15858 hamnavgifter 3
15859 hamnavgifterna 2
15860 hamnbestämmelser 1
15861 hamnen 19
15862 hamninspektioner 1
15863 hamnkategorier 1
15864 hamnkontroll 1
15865 hamnkontrollen 1
15866 hamnmyndigheterna 2
15867 hamnstaten 1
15868 hamra 1
15869 han 1140
15870 hand 147
15871 handbagaget 1
15872 handbojor 1
15873 handdukar 1
15874 handdukarna 1
15875 handel 36
15876 handeln 21
15877 handelns 1
15878 handels- 7
15879 handelsaspekter 1
15880 handelsavtal 9
15881 handelsavtalen 3
15882 handelsavtalet 6
15883 handelsavtalets 1
15884 handelsbalans 1
15885 handelsblockad 1
15886 handelsbolaget 1
15887 handelsfartyg 1
15888 handelsflotta 2
15889 handelsfrågor 3
15890 handelsförbindelser 1
15891 handelsförbindelserna 1
15892 handelsförhandlingar 1
15893 handelsförhandlingarna 1
15894 handelsförmåner 2
15895 handelsglobaliseringen 1
15896 handelshinder 2
15897 handelsintresseaspekten 1
15898 handelsintressen 1
15899 handelskrig 2
15900 handelslogik 1
15901 handelsmässiga 2
15902 handelsmässigt 1
15903 handelsområdet 1
15904 handelsplats 1
15905 handelsplatsen 1
15906 handelsplatser 1
15907 handelspolitik 4
15908 handelspolitiken 2
15909 handelspost 1
15910 handelsreformerna 1
15911 handelsregler 1
15912 handelsreglerna 1
15913 handelsrelaterade 1
15914 handelsrunda 1
15915 handelsrätt 2
15916 handelsrätten 1
15917 handelssamarbete 2
15918 handelssanktioner 1
15919 handelssektorn 1
15920 handelssidan 1
15921 handelssjöfart 1
15922 handelssjöfarten 1
15923 handelsstation 1
15924 handelstvisterna 1
15925 handelsuppgörelser 1
15926 handelsutbyte 4
15927 handelsutbyten 1
15928 handelsutbytespolitik 1
15929 handelsutbytet 3
15930 handelsutveckling 1
15931 handelsvara 4
15932 handelsystem 1
15933 handen 33
15934 handfast 1
15935 handfatet 1
15936 handflata 1
15937 handflatan 1
15938 handflator 1
15939 handfull 4
15940 handha 1
15941 handicap 1
15942 handikapp 8
15943 handikappade 9
15944 handikappades 4
15945 handla 20
15946 handlade 13
15947 handlande 5
15948 handlar 289
15949 handlare 1
15950 handlarna 1
15951 handlas 1
15952 handlat 3
15953 handling 34
15954 handlingar 41
15955 handlingarna 5
15956 handlingen 1
15957 handlingens 1
15958 handlingsalternativ 1
15959 handlingsansvar 1
15960 handlingsfrihet 1
15961 handlingsförlamning 1
15962 handlingsförmåga 3
15963 handlingsförmågan 1
15964 handlingskraft 4
15965 handlingskraftig 1
15966 handlingskraftiga 2
15967 handlingskraftigt 1
15968 handlingslinjer 3
15969 handlingsplan 14
15970 handlingsplanen 4
15971 handlingsplaner 8
15972 handlingsplanernas 1
15973 handlingsprogram 11
15974 handlingsramen 1
15975 handlingssätt 5
15976 handlingssätten 1
15977 handlingssättet 2
15978 handlingsutrymme 5
15979 handläggning 2
15980 handläggningen 2
15981 handpositionerna 1
15982 hands 3
15983 handskarna 1
15984 handskas 13
15985 handske 1
15986 handslaget 1
15987 handtaget 1
15988 handuppräckning 2
15989 handvändning 1
15990 handväska 1
15991 handväskan 1
15992 hankar 1
15993 hans 347
15994 hantera 40
15995 hanterade 1
15996 hanterande 1
15997 hanterandet 1
15998 hanterar 6
15999 hanteras 15
16000 hantering 22
16001 hanteringen 11
16002 hantlangare 1
16003 hantverk 2
16004 hantverkare 2
16005 hantverkarnas 1
16006 hantverksmässiga 2
16007 happy 1
16008 har 5098
16009 haranger 1
16010 haren 1
16011 harmoni 4
16012 harmoniera 1
16013 harmonisera 10
16014 harmoniserad 1
16015 harmoniserade 4
16016 harmoniserar 1
16017 harmoniseras 2
16018 harmoniserat 3
16019 harmoniserats 2
16020 harmonisering 40
16021 harmoniseringen 4
16022 harmoniseringsbegrepp 1
16023 harmoniseringsdirektiv 1
16024 harmonisk 10
16025 harmoniskt 1
16026 harpa 1
16027 hasande 2
16028 hasch 1
16029 hast 2
16030 hastigast 1
16031 hastighet 6
16032 hastigheten 2
16033 hastigheter 2
16034 hastigt 7
16035 hat 2
16036 hatade 1
16037 hatar 1
16038 hatet 3
16039 hatisk 1
16040 hatt 4
16041 hattar 3
16042 hattarna 1
16043 hatten 2
16044 hav 22
16045 havande 1
16046 have 1
16047 have-nots 2
16048 haven 12
16049 havens 2
16050 havererade 1
16051 haveri 5
16052 haveriet 1
16053 haves 2
16054 havet 66
16055 havets 9
16056 havs 23
16057 havs- 1
16058 havsbotten 1
16059 havsdimension 1
16060 havsdäggdjur 1
16061 havsfiske 1
16062 havsforskningsrådet 1
16063 havsföroreningar 2
16064 havsgränsen 1
16065 havsgränser 4
16066 havsgränserna 2
16067 havsinriktning 1
16068 havslivet 1
16069 havsmiljö 4
16070 havsmiljöer 1
16071 havsmiljön 8
16072 havsmiljöns 1
16073 havsnära 1
16074 havsområden 5
16075 havsområdena 1
16076 havsområdenas 1
16077 havsområdet 2
16078 havspolitik 1
16079 havsprodukternas 1
16080 havssköldpaddor 1
16081 havsströmmarna 1
16082 havsvattnet 2
16083 headline 2
16084 hearingen 1
16085 hebreiska 1
16086 heder 2
16087 hederliga 1
16088 hedersamt 1
16089 hederskompani 1
16090 hedersläktaren 1
16091 hedersmedlem 1
16092 hedersplats 1
16093 hedervärt 2
16094 hedga 2
16095 hedniska 1
16096 hedra 5
16097 hedrade 2
16098 hedrande 1
16099 hedrar 1
16100 hejda 2
16101 hejdade 2
16102 hejdas 3
16103 hejdat 1
16104 hejdlösa 1
16105 hektar 3
16106 hektisk 1
16107 hektiska 1
16108 hektometer3 2
16109 hektona 1
16110 hel 43
16111 hela 422
16112 helgar 1
16113 helgdag 1
16114 helgdagar 1
16115 helgedom 1
16116 helgen 2
16117 helgjutna 1
16118 helgon 1
16119 helhet 57
16120 helheten 1
16121 helhetlig 1
16122 helhetsbalansen 1
16123 helhetsbild 2
16124 helhetskoncept 1
16125 helhetslösning 1
16126 helhetspolitik 1
16127 helhetssyn 1
16128 helhetssynen 1
16129 helhjärtad 1
16130 helhjärtade 1
16131 helhjärtat 10
16132 helig 1
16133 heliga 5
16134 helikopter 3
16135 helikoptern 1
16136 helikoptrar 7
16137 helikoptrarna 1
16138 heller 134
16139 hellre 14
16140 hellånga 1
16141 helsike 1
16142 helst 128
16143 helt 415
16144 heltal 1
16145 heltidsanställning 1
16146 heltidsjobb 1
16147 heltäckande 8
16148 heltäckningsmattor 1
16149 helvete 2
16150 helvetesböjda 1
16151 helvetet 1
16152 hem 51
16153 hemarbetet 1
16154 hembygd 1
16155 hemekonomi 1
16156 hemfalla 1
16157 hemförde 1
16158 hemifrån 3
16159 hemkommun 1
16160 hemkänsla 1
16161 hemkära 1
16162 hemland 14
16163 hemlandet 2
16164 hemlig 4
16165 hemliga 7
16166 hemlighet 4
16167 hemligheten 2
16168 hemligheter 3
16169 hemligheterna 1
16170 hemlighetsfulla 1
16171 hemlighetsfullt 3
16172 hemlighålla 2
16173 hemligt 1
16174 hemländer 2
16175 hemläxor 1
16176 hemlösa 7
16177 hemlöshet 3
16178 hemma 23
16179 hemmabasen 1
16180 hemmagjorda 1
16181 hemmamarknad 2
16182 hemmamarknader 2
16183 hemmaplan 1
16184 hemmasittare 1
16185 hemmet 5
16186 hemmets 1
16187 hemort 1
16188 hemregion 2
16189 hemsida 2
16190 hemsk 2
16191 hemska 7
16192 hemskaste 1
16193 hemskickad 1
16194 hemskt 2
16195 hemstad 1
16196 hemställer 1
16197 hemsökelser 1
16198 hemsökt 1
16199 hemvist 2
16200 hemväg 1
16201 henne 87
16202 hennes 101
16203 herodiska 1
16204 heroisk 1
16205 herr 491
16206 herrar 93
16207 herrarna 2
16208 herravälde 2
16209 herraväldet 1
16210 herrelösa 1
16211 herresäte 1
16212 herrgård 1
16213 herrtidningar 1
16214 hertigen 1
16215 hes 2
16216 het 3
16217 heta 6
16218 heter 14
16219 heterogena 1
16220 hets 2
16221 hetsen 1
16222 hett 6
16223 hetta 2
16224 hettan 3
16225 hette 6
16226 hexavalent 1
16227 hibiskus 1
16228 hierarki 1
16229 hierarkin 2
16230 hierarkisering 1
16231 hierarkisk 1
16232 hierarkiska 1
16233 high 3
16234 himlen 10
16235 himmel 5
16236 himmelsskriande 1
16237 hinder 56
16238 hindra 17
16239 hindrade 3
16240 hindrades 1
16241 hindrar 28
16242 hindras 5
16243 hindrat 1
16244 hindrats 1
16245 hindren 3
16246 hindret 1
16247 hinduisk 1
16248 hink 1
16249 hinna 3
16250 hinner 1
16251 hisnande 1
16252 hissade 1
16253 hissen 1
16254 historia 42
16255 historien 18
16256 historiens 3
16257 historier 6
16258 historieskrivningen 1
16259 historik 1
16260 historiker 1
16261 historikern 1
16262 historisk 14
16263 historiska 21
16264 historiskt 12
16265 hit 38
16266 hitintills 1
16267 hitta 61
16268 hittade 8
16269 hittades 2
16270 hittar 13
16271 hittat 6
16272 hittats 1
16273 hittills 98
16274 hittillsvarande 6
16275 hiv-smitta 1
16276 hiv-smittade 1
16277 hivade 1
16278 hjord 2
16279 hjorden 1
16280 hjul 2
16281 hjulen 2
16282 hjulet 1
16283 hjulspår 1
16284 hjälm 1
16285 hjälp 166
16286 hjälpa 104
16287 hjälpande 3
16288 hjälparna 1
16289 hjälpbehov 1
16290 hjälpen 12
16291 hjälper 12
16292 hjälpfunktion 1
16293 hjälpinsatsen 1
16294 hjälpinsatser 3
16295 hjälpkonstruktioner 1
16296 hjälplösa 2
16297 hjälplöst 2
16298 hjälpmedel 2
16299 hjälporganisationer 1
16300 hjälpprogram 1
16301 hjälpt 3
16302 hjälpta 1
16303 hjälpte 4
16304 hjälptjänster 1
16305 hjälpvilliga 1
16306 hjältar 4
16307 hjälten 1
16308 hjärna 1
16309 hjärnkapacitet 1
16310 hjärnor 2
16311 hjärnorna 1
16312 hjärta 8
16313 hjärtan 4
16314 hjärtans 3
16315 hjärtat 15
16316 hjärtliga 2
16317 hjärtligt 19
16318 hjärtpunkt 1
16319 hjärtstoppande 1
16320 hjässa 2
16321 hoande 1
16322 hobby 2
16323 hobbybilar 1
16324 hoc-direktiv 1
16325 hoc-transporter 1
16326 hojtade 1
16327 holländsk 1
16328 holländska 2
16329 home 1
16330 homofobin 1
16331 homogen 1
16332 homogena 1
16333 homogent 4
16334 homosexuell 1
16335 homosexuella 1
16336 hon 267
16337 honnör 1
16338 honom 305
16339 hop 1
16340 hopas 1
16341 hope 1
16342 hopfällbart 1
16343 hopkok 1
16344 hopp 22
16345 hoppa 2
16346 hoppade 5
16347 hoppades 7
16348 hoppar 1
16349 hoppas 286
16350 hoppats 2
16351 hoppet 5
16352 hoppfullhet 1
16353 hoppingivande 3
16354 hopplös 1
16355 hopplöst 6
16356 hora 1
16357 hord 1
16358 horderna 1
16359 horisont 1
16360 horisontala 2
16361 horisontella 4
16362 horisontellt 3
16363 horisonten 3
16364 hormonbehandlat 1
16365 hormonstörande 2
16366 horn 2
16367 hornen 1
16368 hos 194
16369 hospice 1
16370 hostade 2
16371 hot 31
16372 hota 2
16373 hotad 4
16374 hotade 6
16375 hotades 3
16376 hotande 4
16377 hotar 25
16378 hotas 15
16379 hotat 2
16380 hotats 2
16381 hotbilden 1
16382 hotbilder 1
16383 hotell 1
16384 hotell- 1
16385 hotellen 1
16386 hotellet 3
16387 hotellets 1
16388 hotellägare 1
16389 hotelser 2
16390 hotet 10
16391 hotfull 1
16392 hotfulla 1
16393 hotfullt 1
16394 http://officeupdate.microsoft.com/ 1
16395 hud 1
16396 huden 2
16397 hudfärg 3
16398 hugg 3
16399 hugga 1
16400 huggas 1
16401 hukade 3
16402 huliganerna 1
16403 human 2
16404 humanism 1
16405 humanistiska 2
16406 humanitet 1
16407 humanitär 14
16408 humanitära 19
16409 humanitäras 2
16410 humanitärt 4
16411 humankapital 3
16412 humankapitalet 1
16413 humbug 1
16414 humlen 1
16415 humor 1
16416 humör 2
16417 hund 4
16418 hundar 1
16419 hundbajs 1
16420 hunden 2
16421 hundens 1
16422 hundra 10
16423 hundrade 1
16424 hundrafemtio 1
16425 hundraprocentig 2
16426 hundraprocentigt 1
16427 hundraser 1
16428 hundratal 1
16429 hundratals 12
16430 hundratusentals 12
16431 hundskall 1
16432 hunger 2
16433 hungersnöd 2
16434 hungrig 3
16435 hungrigare 1
16436 hunnit 4
16437 hur 558
16438 hurdan 2
16439 huruvida 27
16440 hus 32
16441 husalf 2
16442 husalfer 1
16443 husarrest 1
16444 husbonde 1
16445 husdjur 1
16446 husen 2
16447 huset 22
16448 husets 3
16449 hushåll 5
16450 hushålla 1
16451 hushållen 1
16452 hushållning 2
16453 hushålls- 1
16454 hushållsvatten 1
16455 hushållsändamål 1
16456 husligt 1
16457 husrum 1
16458 hustak 1
16459 hustru 16
16460 hustrun 4
16461 hustruns 1
16462 husövertaganden 1
16463 huva 1
16464 huvan 1
16465 huvud 48
16466 huvudaktiviteter 1
16467 huvudaktör 1
16468 huvudangelägenheter 1
16469 huvudansvaret 5
16470 huvudargument 1
16471 huvudbeståndsdelar 1
16472 huvudbudskap 2
16473 huvudbyggnad 1
16474 huvudbyggnaden 1
16475 huvuddel 1
16476 huvuddelen 1
16477 huvuddrag 1
16478 huvuddragen 3
16479 huvuden 4
16480 huvudena 1
16481 huvudet 22
16482 huvudfinansieringen 1
16483 huvudfråga 4
16484 huvudfrågan 1
16485 huvudförslagen 1
16486 huvudinriktning 1
16487 huvudinriktningar 1
16488 huvudkontor 3
16489 huvudkravet 1
16490 huvudlinjerna 2
16491 huvudmål 3
16492 huvudpersonerna 1
16493 huvudprincip 1
16494 huvudpunkter 1
16495 huvudrekommendationer 1
16496 huvudroll 3
16497 huvudrollsinnehavarna 1
16498 huvudrubriker 1
16499 huvudrätten 1
16500 huvudsak 18
16501 huvudsaken 2
16502 huvudsakliga 15
16503 huvudsaklige 1
16504 huvudsakligen 30
16505 huvudskälet 1
16506 huvudstad 4
16507 huvudstaden 3
16508 huvudstadens 1
16509 huvudstäder 2
16510 huvudstäderna 3
16511 huvudsyfte 1
16512 huvudsyften 1
16513 huvudsyftet 1
16514 huvudtaget 1
16515 huvuduppgift 1
16516 huvuduppgifter 1
16517 huvudvärk 2
16518 hy 5
16519 hybridbetänkande 1
16520 hycklade 1
16521 hycklande 4
16522 hyckleri 8
16523 hyckleriet 2
16524 hydda 1
16525 hyddan 1
16526 hyddor 2
16527 hydrauliska 1
16528 hydrogeologiskt 1
16529 hydrologiska 1
16530 hygglig 1
16531 hygien 3
16532 hygienens 1
16533 hygieniska 1
16534 hylla 5
16535 hyllade 1
16536 hyllan 1
16537 hyllandet 1
16538 hyllar 1
16539 hyllas 1
16540 hyllning 2
16541 hylsa 1
16542 hypereffektiva 1
16543 hyperlänkarna 1
16544 hypnotiserade 2
16545 hypotes 1
16546 hypotesen 1
16547 hypoteser 1
16548 hypotetiska 1
16549 hypotetiskt 2
16550 hyr 1
16551 hyrd 1
16552 hyreshus 1
16553 hysa 7
16554 hyser 10
16555 hyste 1
16556 hysterin 1
16557 hytt 1
16558 hytten 2
16559 häck 1
16560 häcken 7
16561 hädanefter 2
16562 hädelser 2
16563 häftiga 4
16564 häftigt 2
16565 hägn 1
16566 häktade 1
16567 häktningen 1
16568 häktningsorder 1
16569 häl 2
16570 häleri 1
16571 hälft 2
16572 hälften 19
16573 hällde 2
16574 hälsa 50
16575 hälsade 7
16576 hälsades 2
16577 hälsan 8
16578 hälsar 9
16579 hälsning 1
16580 hälsningar 2
16581 hälsningen 1
16582 hälso- 6
16583 hälsoaspekten 1
16584 hälsobehoven 1
16585 hälsobringande 1
16586 hälsoeffekter 1
16587 hälsoeffekterna 1
16588 hälsofrämjande 1
16589 hälsofrågor 3
16590 hälsoområden 1
16591 hälsoproblem 1
16592 hälsoproblemen 1
16593 hälsorelaterade 1
16594 hälsorisker 1
16595 hälsosam 2
16596 hälsosamma 1
16597 hälsosektorn 3
16598 hälsosituationen 1
16599 hälsoskydd 3
16600 hälsoskyddet 1
16601 hälsosystemet 1
16602 hälsotillstånd 3
16603 hälsotjänster 1
16604 hälsovådliga 1
16605 hälsovård 13
16606 hälsovården 3
16607 hälsovårdsanordningar 1
16608 hälsovårdsdepartement 1
16609 hälsovårdsinrättningar 2
16610 hälsovårdsinspektören 1
16611 hälsovårdskostnader 1
16612 hälsovårdsområdet 1
16613 hälsovårdssystem 2
16614 hälsovårdssystemet 3
16615 hämma 1
16616 hämmar 2
16617 hämmas 1
16618 hämnande 1
16619 hämnas 2
16620 hämnd 2
16621 hämndbegär 1
16622 hämndlystnad 1
16623 hämningslös 1
16624 hämta 11
16625 hämtad 1
16626 hämtade 2
16627 hämtar 2
16628 hämtas 4
16629 hämtat 2
16630 hämtning 1
16631 hända 34
16632 hände 33
16633 händelse 31
16634 händelseförloppet 1
16635 händelselös 1
16636 händelsemönster 1
16637 händelsen 7
16638 händelsens 1
16639 händelser 39
16640 händelserikt 1
16641 händelserna 17
16642 händelseutveckling 1
16643 händelseutvecklingen 1
16644 händelsevis 2
16645 händer 61
16646 händerna 23
16647 händigt 1
16648 hänför 2
16649 hänförde 1
16650 hänga 5
16651 hängande 4
16652 hängbro 1
16653 hängde 17
16654 hänge 3
16655 hänger 28
16656 hängett 1
16657 hängivelse 1
16658 hängivenhet 1
16659 hänglås 1
16660 hängning 1
16661 hängslen 1
16662 hänseende 15
16663 hänseenden 4
16664 hänseendet 4
16665 hänskjuta 1
16666 hänsyn 200
16667 hänsynen 5
16668 hänsynsfull 1
16669 hänsynslös 1
16670 hänsynstaganden 3
16671 hänsynstagandet 3
16672 hänt 27
16673 hänvisa 20
16674 hänvisad 1
16675 hänvisade 18
16676 hänvisades 2
16677 hänvisar 22
16678 hänvisas 5
16679 hänvisat 6
16680 hänvisats 3
16681 hänvisning 25
16682 hänvisningar 8
16683 hänvisningarna 1
16684 hänvisningen 8
16685 häpen 1
16686 häpnad 3
16687 häpnadsväckande 1
16688 häpnar 1
16689 här 1145
16690 härden 1
16691 härefter 1
16692 häri 1
16693 härifrån 3
16694 härigenom 4
16695 härjade 2
16696 härledas 2
16697 härliga 1
16698 härligaste 1
16699 härligt 1
16700 härmade 2
16701 härmed 12
16702 häromdagen 1
16703 härrör 19
16704 härs 1
16705 härskar 1
16706 härskare 2
16707 härskarinnan 1
16708 härskarna 1
16709 härskaror 1
16710 härstammar 7
16711 härtill 1
16712 härutöver 1
16713 härva 1
16714 härvidlag 1
16715 häst 5
16716 hästar 2
16717 hästen 4
16718 hästkapplöpning 1
16719 hästliknande 1
16720 hästskor 1
16721 häva 5
16722 hävas 3
16723 hävda 18
16724 hävdade 8
16725 hävdar 22
16726 hävdas 1
16727 hävdat 7
16728 hävdvunna 1
16729 häver 2
16730 hävning 1
16731 hävstången 1
16732 hävts 1
16733 häxa 3
16734 häxan 1
16735 häxkonst 1
16736 häxkonster 1
16737 häxor 2
16738 hågen 1
16739 håglöst 1
16740 hål 5
16741 håla 1
16742 håll 48
16743 hålla 101
16744 hållas 14
16745 hållbar 85
16746 hållbara 15
16747 hållbarhet 5
16748 hållbart 18
16749 hållen 2
16750 håller 190
16751 hållet 39
16752 hållit 18
16753 hållits 3
16754 hållna 2
16755 hållning 24
16756 hållningen 2
16757 hållplats 1
16758 hålls 14
16759 hålor 1
16760 hån 2
16761 hånade 1
16762 hånar 1
16763 hånflinande 1
16764 hånfull 1
16765 hånglat 1
16766 hår 22
16767 hård 13
16768 hårda 16
16769 hårdare 5
16770 hårdast 4
16771 hårdhandskarna 1
16772 hårdingar 1
16773 hårdingen 1
16774 hårdnackade 1
16775 hårdnackat 2
16776 hårdvara 1
16777 håret 12
16778 hårfina 1
16779 hårklyverier 1
16780 hårnät 1
16781 hårnål 1
16782 hårnålar 1
16783 hårnålen 1
16784 hårstrå 2
16785 hårt 48
16786 hårtestar 1
16787 håvar 1
16788 höft 1
16789 höfterna 1
16790 hög 106
16791 höga 65
16792 högaktar 1
16793 högaktuellt 1
16794 högar 1
16795 höge 34
16796 höger 13
16797 högerextremismen 1
16798 högerextremismens 1
16799 högerextremistiska 3
16800 högerhanden 1
16801 högerkanten 1
16802 högerkvinnor 1
16803 högerledamöters 1
16804 högermajoritet 1
16805 högern 5
16806 högerns 4
16807 högerpopulists 1
16808 högervridning 1
16809 högg 1
16810 höghastighetståg 1
16811 höginkomstländer 1
16812 höginkomsttagare 1
16813 högkonjunktur 1
16814 högkostnadsområden 1
16815 högkvalitativ 2
16816 högkvalitativa 1
16817 högkvarter 1
16818 högljudd 1
16819 högljudda 1
16820 högljutt 2
16821 högländerna 2
16822 högnivågrupp 3
16823 högnivågruppen 6
16824 högprestationstjänst 1
16825 högpresterande 1
16826 högra 2
16827 högre 78
16828 högrest 1
16829 högriskfonder 1
16830 högriskprodukter 1
16831 högröda 1
16832 högrörliga 1
16833 högskolor 1
16834 högst 37
16835 högsta 38
16836 högste 1
16837 högstämda 1
16838 högstärkelsekrage 1
16839 högt 40
16840 högteknologiska 2
16841 högtidliga 1
16842 högtidligen 1
16843 högtidligheten 1
16844 högtidlighålla 1
16845 högtidligt 8
16846 högtravande 2
16847 höja 15
16848 höjas 5
16849 höjd 8
16850 höjda 2
16851 höjde 2
16852 höjden 2
16853 höjderna 1
16854 höjdpunkt 2
16855 höjdpunkten 1
16856 höjer 3
16857 höjning 7
16858 höjningar 1
16859 höjningen 3
16860 höjs 2
16861 höjt 1
16862 höjts 1
16863 hölje 1
16864 höljs 1
16865 höll 47
16866 hölls 8
16867 höna 1
16868 hönor 1
16869 hör 92
16870 höra 71
16871 hörande 1
16872 höras 5
16873 hörbar 1
16874 hörbart 1
16875 hörd 4
16876 hörda 1
16877 hörde 37
16878 hördes 11
16879 hörn 6
16880 hörnen 2
16881 hörnet 5
16882 hörnsten 2
16883 hörnstenen 1
16884 hörsammar 1
16885 hörsammats 2
16886 hört 76
16887 hörts 3
16888 höst 2
16889 höstack 1
16890 höstas 2
16891 hösten 3
16892 hövlig 1
16893 hövlighet 1
16894 i 12839
16895 i- 1
16896 iaktta 10
16897 iakttagande 4
16898 iakttagelse 1
16899 iakttagelser 4
16900 iakttagelserna 1
16901 iakttagit 1
16902 iakttar 2
16903 iakttas 6
16904 iakttog 3
16905 ianspråktagandet 1
16906 iberiska 1
16907 ibland 65
16908 icke 41
16909 icke- 1
16910 icke-albaner 1
16911 icke-albanska 3
16912 icke-avvisning 1
16913 icke-bergsregioner 1
16914 icke-budgetisering 1
16915 icke-danska 1
16916 icke-diskriminerande 1
16917 icke-diskriminering 3
16918 icke-dokument 1
16919 icke-européer- 1
16920 icke-fossil 1
16921 icke-handikappade 1
16922 icke-harmoniserade 3
16923 icke-inblandning 1
16924 icke-införlivande 1
16925 icke-insatta 1
16926 icke-intervention 1
16927 icke-interventionsmotionen 1
16928 icke-kommersiella 1
16929 icke-kvalificerade 1
16930 icke-lönerelaterade 1
16931 icke-magiska 1
16932 icke-medborgare 1
16933 icke-medlemsstater 1
16934 icke-metalldelar 1
16935 icke-militära 1
16936 icke-rasistiskt 1
16937 icke-regeringssektorns 1
16938 icke-självvalda 1
16939 icke-spridningsavtalet 3
16940 icke-statlig 1
16941 icke-statliga 40
16942 icke-statligt 1
16943 icke-tariffiära 1
16944 icke-tillämpning 1
16945 icke-ömsesidiga 1
16946 ickenylonhud 1
16947 ickesjälsligt 1
16948 idag 12
16949 ideal 4
16950 ideala 2
16951 idealen 2
16952 idealet 2
16953 idealiserat 1
16954 idealisk 1
16955 idealiska 1
16956 idealiskt 1
16957 idealism 2
16958 idealistiskt 1
16959 ideella 2
16960 idel 1
16961 ideligen 2
16962 identifiera 13
16963 identifierade 4
16964 identifierades 1
16965 identifierar 5
16966 identifieras 4
16967 identifierat 7
16968 identifierats 1
16969 identifierbara 1
16970 identifiering 1
16971 identifieringen 1
16972 identifikation 1
16973 identisk 1
16974 identiska 1
16975 identiskt 1
16976 identitet 16
16977 identiteten 3
16978 identiteter 3
16979 identitetshandlingar 2
16980 ideolog 1
16981 ideologi 4
16982 ideologisk 2
16983 ideologiska 7
16984 ideologiskt 2
16985 idiosynkrasi 1
16986 idiot 4
16987 idioterna 1
16988 idiotisk 1
16989 idiotiska 1
16990 idrott 5
16991 idrottssammanhang 1
16992 idyllisk 1
16993 idé 27
16994 idéer 35
16995 idéerna 1
16996 idén 32
16997 ifall 7
16998 ifråga 3
16999 ifrågasatt 1
17000 ifrågasatte 1
17001 ifrågasattes 2
17002 ifrågasatts 1
17003 ifrågasätta 13
17004 ifrågasättande 3
17005 ifrågasättanden 1
17006 ifrågasättandet 1
17007 ifrågasättas 4
17008 ifrågasätter 12
17009 ifrågasätts 7
17010 ifrågavarande 4
17011 ifrån 74
17012 iförd 4
17013 igelkott 1
17014 igen 146
17015 igenkännande 3
17016 igenom 69
17017 igenom- 1
17018 igenspikade 1
17019 ignorera 4
17020 ignorerade 2
17021 ignorerades 1
17022 ignoreras 3
17023 igång 29
17024 igångkörning 1
17025 igångsättandet 2
17026 igår 1
17027 ihjäl 3
17028 ihop 49
17029 ihopsatt 1
17030 ihärdighet 1
17031 ihåg 49
17032 ihåliga 1
17033 ihållande 8
17034 ikapp 1
17035 ikraftträdande 4
17036 ikraftträdandet 3
17037 ikväll 1
17038 il 1
17039 illa 19
17040 illaluktande 1
17041 illavarslande 2
17042 illegal 5
17043 illegala 12
17044 illegalt 5
17045 illojal 1
17046 illojala 2
17047 illusion 4
17048 illusionen 1
17049 illusioner 1
17050 illusionism 1
17051 illusionsfrie 1
17052 illusoriskt 1
17053 illustration 2
17054 illustrera 3
17055 illustrerade 1
17056 illustrerar 1
17057 illustreras 2
17058 illvilliga 1
17059 illvilligt 2
17060 ilska 4
17061 ilsken 1
17062 ilsket 3
17063 ilskna 2
17064 image 1
17065 imaginära 1
17066 imitationsprodukter 1
17067 imitera 1
17068 immaterialrätt 3
17069 immaterialrätten 3
17070 immaterialrättsliga 2
17071 immaterialrättsligt 2
17072 immateriella 5
17073 immigrantbefolkningen 1
17074 immigranter 3
17075 immigration 3
17076 immigrationen 1
17077 immigrationsblanketterna 1
17078 immigrationspolitiken 1
17079 immigrationsprocess 1
17080 immunitet 7
17081 immuniteten 5
17082 imperativ 2
17083 imperialisternas 1
17084 imperialistiska 1
17085 imperiebyggare 1
17086 implementation 1
17087 implementerade 2
17088 implementeringen 2
17089 implicit 1
17090 impolitiskt 1
17091 imponera 1
17092 imponerad 1
17093 imponerade 1
17094 imponerande 3
17095 impopulära 1
17096 impopulärt 1
17097 import 6
17098 importbegränsningarna 1
17099 importen 5
17100 importera 8
17101 importerad 3
17102 importerade 3
17103 importerar 2
17104 importeras 5
17105 importerats 1
17106 importförbudet 1
17107 importhinder 1
17108 importpolitik 2
17109 importrestriktioner 1
17110 importsystemet 1
17111 impossible 1
17112 improviserat 1
17113 impuls 4
17114 impulsen 1
17115 impulser 11
17116 impulsiv 1
17117 impunity 1
17118 in 436
17119 in- 1
17120 inaktiverat 1
17121 inaktivt 1
17122 inarbetats 1
17123 inbegripa 6
17124 inbegripande 1
17125 inbegripandet 1
17126 inbegripas 3
17127 inbegripen 1
17128 inbegriper 18
17129 inbegripet 20
17130 inbegripna 2
17131 inbegrips 2
17132 inbesparingar 1
17133 inbilla 2
17134 inbillad 1
17135 inbillade 1
17136 inbjuda 2
17137 inbjudan 2
17138 inbjudande 1
17139 inbjuden 2
17140 inbjuder 3
17141 inbjudit 1
17142 inbjudits 1
17143 inbjudna 2
17144 inbjudningar 1
17145 inbjöd 1
17146 inblandad 3
17147 inblandade 20
17148 inblandat 3
17149 inblandning 22
17150 inbringade 2
17151 inbringar 1
17152 inbyggd 2
17153 inbyggt 1
17154 inbördes 21
17155 inbördeskrig 3
17156 inbördeskriget 3
17157 incheckningstid 1
17158 incident 1
17159 incitament 14
17160 incitamenten 2
17161 incitamentet 4
17162 indelade 2
17163 indelas 2
17164 indelat 1
17165 index 2
17166 indexering 2
17167 indexet 1
17168 indexfond 1
17169 indianer 1
17170 indianerna 2
17171 indianernas 1
17172 indianska 1
17173 indicier 2
17174 indignation 3
17175 indignerad 1
17176 indikation 1
17177 indikationer 1
17178 indikativt 1
17179 indikatorer 12
17180 indikatorn 1
17181 indirekt 15
17182 indirekta 6
17183 indiska 2
17184 indiskret 1
17185 individ 7
17186 individen 1
17187 individens 3
17188 individer 10
17189 individerna 1
17190 individers 1
17191 individs 1
17192 individualiserade 1
17193 individualisering 1
17194 individualism 2
17195 individualitet 1
17196 individuell 2
17197 individuella 14
17198 individuellt 2
17199 indonesisk 1
17200 indonesiska 1
17201 indonesiskt 1
17202 indraget 1
17203 indragning 1
17204 indränkt 1
17205 industri 16
17206 industri- 4
17207 industrial 1
17208 industrialiserade 2
17209 industrialiseringen 1
17210 industriell 2
17211 industriella 11
17212 industriellt 1
17213 industrier 7
17214 industrierna 1
17215 industriernas 1
17216 industrifrågor 6
17217 industriföretagen 1
17218 industriföroreningar 1
17219 industrigrupper 1
17220 industrikatastrofer 1
17221 industrikulturen 1
17222 industriliknande 1
17223 industrilobbyisten 1
17224 industriländerna 2
17225 industrimässor 1
17226 industrin 38
17227 industrins 4
17228 industripolitikerna 1
17229 industripolitisk 1
17230 industriprodukt 1
17231 industriprodukter 1
17232 industris 1
17233 industrisektorer 1
17234 industriverksamheten 1
17235 industriverksamheter 1
17236 indämda 1
17237 ineffektiv 2
17238 ineffektiva 5
17239 ineffektivitet 4
17240 ineffektivt 2
17241 infallsvinklar 1
17242 infallsvinklarna 1
17243 infann 1
17244 infantiliserande 1
17245 infekterade 2
17246 infektion 1
17247 infektionsnivåer 1
17248 infektionssjukdom 1
17249 infektiös 5
17250 infernaliska 2
17251 inferno 2
17252 infernos 1
17253 infiltrera 1
17254 infinitum 1
17255 infinner 1
17256 inflation 6
17257 inflationen 8
17258 inflationsbekämpning 1
17259 inflationsbekämpningen 1
17260 inflationstakten 1
17261 inflationstrycket 1
17262 influerad 1
17263 inflytande 24
17264 inflytelserika 1
17265 infogas 1
17266 information 153
17267 informationen 39
17268 informationer 1
17269 informations- 13
17270 informationsanalys 1
17271 informationsanalytiker 1
17272 informationsbrist 1
17273 informationsbudget 2
17274 informationsbärare 1
17275 informationscentrerna 1
17276 informationscentrum 1
17277 informationsekonomi 1
17278 informationsfattiga 1
17279 informationsflöde 1
17280 informationsfrihet 2
17281 informationsfrågan 1
17282 informationsinsamling 2
17283 informationskampanj 4
17284 informationskampanjen 2
17285 informationskampanjer 1
17286 informationskanal 1
17287 informationsmöte 1
17288 informationspolitik 1
17289 informationspolitiken 1
17290 informationsproblem 1
17291 informationsrika 1
17292 informationssamhälle 2
17293 informationssamhället 16
17294 informationssamhällets 1
17295 informationssystem 7
17296 informationsteknik 6
17297 informationstekniken 6
17298 informationsteknikmarknaderna 1
17299 informationsteknisk 1
17300 informationstekniska 2
17301 informationsteknologi 1
17302 informationsteknologin 4
17303 informationsutbyte 5
17304 informationsutbytet 4
17305 informationsvilja 1
17306 informationsåtgärder 2
17307 informationsöverföringens 1
17308 informella 7
17309 informellt 2
17310 informera 30
17311 informerad 3
17312 informerade 10
17313 informerades 2
17314 informerar 1
17315 informeras 6
17316 informerat 5
17317 informerats 3
17318 infrastruktur 22
17319 infrastrukturbestämmelser 1
17320 infrastrukturell 1
17321 infrastrukturella 1
17322 infrastrukturen 7
17323 infrastrukturens 2
17324 infrastrukturer 11
17325 infrastrukturerna 2
17326 infrastrukturnätet 1
17327 infrastrukturprogram 1
17328 infrastrukturprojekt 1
17329 infrastruktursatsningar 1
17330 infrastrukturutvecklingen 1
17331 infrastrukturåtgärder 1
17332 infria 1
17333 infriade 1
17334 infriades 1
17335 infrias 1
17336 infunnit 2
17337 infällda 1
17338 infångad 1
17339 infödda 1
17340 infödingarna 2
17341 inföll 1
17342 inför 279
17343 införa 96
17344 införande 8
17345 införandet 24
17346 införas 18
17347 införde 3
17348 infördes 5
17349 införliva 16
17350 införlivade 1
17351 införlivades 4
17352 införlivande 11
17353 införlivandet 9
17354 införlivar 3
17355 införlivas 15
17356 införlivat 1
17357 införlivats 5
17358 införs 9
17359 införsel 2
17360 införselrestriktioner 1
17361 införstådd 2
17362 införstådda 1
17363 infört 11
17364 införts 7
17365 inga 101
17366 ingalunda 6
17367 ingav 2
17368 ingavs 2
17369 inge 2
17370 ingefära 1
17371 ingen 228
17372 ingenjör 2
17373 ingenjörer 1
17374 ingenstans 5
17375 ingenting 92
17376 inger 6
17377 inget 98
17378 ingett 2
17379 ingick 3
17380 ingivit 8
17381 ingivits 3
17382 ingjuta 1
17383 ingrediens 1
17384 ingredienser 3
17385 ingrep 1
17386 ingrepp 9
17387 ingreppen 2
17388 ingress 1
17389 ingressen 1
17390 ingripa 20
17391 ingripande 13
17392 ingripanden 1
17393 ingripandet 1
17394 ingriper 3
17395 ingripit 4
17396 ingrott 1
17397 ingå 24
17398 ingående 15
17399 ingångar 1
17400 ingår 49
17401 ingått 8
17402 ingåtts 4
17403 inhemsk 1
17404 inhemska 12
17405 inhämta 2
17406 inhämtande 1
17407 inhämtar 1
17408 inhämtas 1
17409 inhämtat 1
17410 inifrån 4
17411 initiativ 161
17412 initiativandan 1
17413 initiativbetänkande 2
17414 initiativen 7
17415 initiativet 35
17416 initiativets 1
17417 initiativförmåga 1
17418 initiativkraft 2
17419 initiativrik 1
17420 initiativrikt 1
17421 initiativrätt 8
17422 initiativrätten 2
17423 initiativs 1
17424 initiativtagares 1
17425 initiera 1
17426 initierade 1
17427 initierades 1
17428 initierat 3
17429 injicerats 1
17430 inkapslade 2
17431 inkarnationen 2
17432 inkilade 1
17433 inkludera 12
17434 inkluderade 1
17435 inkluderades 1
17436 inkluderandet 1
17437 inkluderar 5
17438 inkluderas 5
17439 inkluderat 3
17440 inkluderats 1
17441 inklusive 49
17442 inkom 1
17443 inkompetens 3
17444 inkompetensen 1
17445 inkompetenta 1
17446 inkomst 7
17447 inkomst- 1
17448 inkomsten 2
17449 inkomster 17
17450 inkomsterna 3
17451 inkomstfördelning 1
17452 inkomstförluster 1
17453 inkomstkälla 4
17454 inkomstkällor 1
17455 inkomstskapande 1
17456 inkomststöd 1
17457 inkonsekvens 1
17458 inkonsekvenser 1
17459 inkonsekvenserna 1
17460 inkonsekvent 1
17461 inkorporera 1
17462 inkorrekta 1
17463 inkräkta 1
17464 inkubationsperiod 1
17465 inköp 3
17466 inköpsbesluten 1
17467 inköpslistor 2
17468 inköpslistorna 1
17469 inkörsport 1
17470 inlandet 1
17471 inlands- 1
17472 inlandsstaterna 1
17473 inleda 61
17474 inledande 8
17475 inledandet 2
17476 inledas 9
17477 inledde 9
17478 inleddes 11
17479 inleder 12
17480 inledning 2
17481 inledningen 10
17482 inledningsanförande 1
17483 inledningsfasen 1
17484 inledningsskedet 3
17485 inledningsvis 8
17486 inleds 12
17487 inlett 10
17488 inletts 20
17489 inloggningskonton 1
17490 inloggningslösenord 1
17491 inloggningsnamn 1
17492 inlägg 42
17493 inlägga 1
17494 inläggen 4
17495 inlägget 2
17496 inlämnade 2
17497 inlämnades 2
17498 inlämnande 1
17499 inlämning 3
17500 inlämnings- 1
17501 inlämningsdatumen 1
17502 inlärningsproblem 1
17503 inlåst 1
17504 inlåsta 1
17505 inlåta 1
17506 inlåter 1
17507 inlöpande 1
17508 innan 135
17509 innandömen 2
17510 innanför 7
17511 inne 25
17512 inne-semantik 1
17513 innebar 8
17514 inneboende 3
17515 inneburit 3
17516 innebär 257
17517 innebära 59
17518 innebörd 4
17519 innebörden 12
17520 innefatta 1
17521 innefattade 1
17522 innefattande 1
17523 innefattar 12
17524 innefattas 8
17525 innehaft 1
17526 innehar 12
17527 innehas 2
17528 innehav 1
17529 innehavarna 1
17530 innehavet 1
17531 innehåll 32
17532 innehålla 19
17533 innehållande 2
17534 innehåller 100
17535 innehållet 51
17536 innehållit 2
17537 innehållsdeklaration 1
17538 innehållsindustrin 1
17539 innehållslig 1
17540 innehållsliga 3
17541 innehållsmässigt 2
17542 innehållsrika 2
17543 innehöll 10
17544 inneperiod 1
17545 innerfickan 1
17546 innerliga 3
17547 innerligt 3
17548 innerst 1
17549 innersta 2
17550 innerstad 1
17551 innersulor 1
17552 innevarande 3
17553 innevånare 2
17554 innovation 16
17555 innovationer 4
17556 innovationsföretag 1
17557 innovationspolitik 1
17558 innovationsprojekt 1
17559 innovativ 5
17560 innovativa 14
17561 innovativt 1
17562 innovatörer 1
17563 innovatörerna 1
17564 inofficiella 1
17565 inom 894
17566 inombords 2
17567 inomeuropeiska 1
17568 inomhustoalett 1
17569 inpränta 1
17570 inpräntat 1
17571 inpå 2
17572 inramad 1
17573 inramade 2
17574 inramning 2
17575 inre 203
17576 inresa 3
17577 inrikes 21
17578 inrikes- 3
17579 inrikesfrågor 2
17580 inrikesminister 1
17581 inrikesministeriet 1
17582 inrikesministern 3
17583 inrikesministrar 1
17584 inrikesministrarna 1
17585 inrikespolitik 3
17586 inrikespolitiska 3
17587 inrikta 14
17588 inriktad 10
17589 inriktade 5
17590 inriktar 5
17591 inriktas 5
17592 inriktat 5
17593 inriktning 32
17594 inriktningar 5
17595 inriktningen 10
17596 inrotad 1
17597 inryms 2
17598 inrätta 54
17599 inrättade 4
17600 inrättades 6
17601 inrättande 5
17602 inrättandet 22
17603 inrättar 6
17604 inrättas 13
17605 inrättat 3
17606 inrättats 5
17607 inrättningar 4
17608 inrättningarna 2
17609 inrådan 1
17610 insamlade 2
17611 insamlas 2
17612 insamling 19
17613 insamlingen 2
17614 insamlingsanläggning 1
17615 insamlingsmetoderna 1
17616 insats 36
17617 insatsen 3
17618 insatser 75
17619 insatserna 20
17620 insatsområden 1
17621 insatsområdena 1
17622 insatsstyrka 3
17623 insatsstyrkan 4
17624 insatt 1
17625 inse 32
17626 insegel 1
17627 insekter 2
17628 insektsmedel 1
17629 inser 41
17630 insett 4
17631 insikt 4
17632 insikten 4
17633 insikter 1
17634 insiktsfulla 1
17635 insistera 17
17636 insisterade 2
17637 insisterar 10
17638 inskickandet 1
17639 inskrida 1
17640 inskriven 2
17641 inskränka 6
17642 inskränkande 1
17643 inskränker 7
17644 inskränkning 3
17645 inskränkningar 4
17646 inskränkningarna 2
17647 inskränks 1
17648 inskränkte 1
17649 inskränkts 1
17650 inslag 11
17651 inslagen 3
17652 inslaget 2
17653 inslagna 2
17654 insläppningsknappen 1
17655 insnärjda 1
17656 insolvens 4
17657 insolvensförfarande 1
17658 insolvensförfaranden 2
17659 inspekterades 1
17660 inspekteras 1
17661 inspektion 2
17662 inspektioner 4
17663 inspektionerna 1
17664 inspektionsmyndigheterna 1
17665 inspektionssystem 1
17666 inspektörer 5
17667 inspektörernas 1
17668 inspektörskår 1
17669 inspiration 1
17670 inspirationskällor 1
17671 inspiratörer 1
17672 inspirerad 1
17673 inspirerande 1
17674 inspireras 1
17675 inspirerat 1
17676 inspirerats 1
17677 inspärrade 1
17678 instabil 3
17679 instabila 1
17680 instabilitet 3
17681 instabiliteten 1
17682 installationerna 1
17683 installationsalternativ 1
17684 installationssidan 1
17685 installera 4
17686 installerade 2
17687 installeras 4
17688 installerat 5
17689 installerats 2
17690 instans 5
17691 instanser 9
17692 instanserna 7
17693 insteg 1
17694 instifta 2
17695 instiftats 1
17696 instinkt 1
17697 instinkter 1
17698 instinktiva 1
17699 instituten 2
17700 institution 28
17701 institutionell 9
17702 institutionella 32
17703 institutionellt 3
17704 institutionen 3
17705 institutionens 1
17706 institutioner 94
17707 institutionerna 76
17708 institutionernas 12
17709 institutioners 7
17710 institutionsansvariga 1
17711 institutionsprojekt 1
17712 institutionsreformen 1
17713 instruktioner 2
17714 instrument 110
17715 instrumentaliseras 1
17716 instrumentbrädan 1
17717 instrumenten 10
17718 instrumenterad 1
17719 instrumentet 15
17720 instrumentets 1
17721 instruments 2
17722 inställa 4
17723 inställd 9
17724 inställda 4
17725 inställer 3
17726 inställning 55
17727 inställningar 1
17728 inställningarna 1
17729 inställningen 12
17730 inställsamma 1
17731 inställsamt 2
17732 inställt 2
17733 instämde 2
17734 instämma 13
17735 instämmande 4
17736 instämmer 41
17737 instängd 1
17738 instängda 2
17739 instängt 1
17740 insvept 1
17741 insyn 23
17742 insynen 3
17743 insynsskyddat 1
17744 insändare 1
17745 insättande 1
17746 insättningar 1
17747 insåg 12
17748 inta 15
17749 intagit 6
17750 intagits 1
17751 intakta 1
17752 intala 1
17753 intar 13
17754 intas 2
17755 inte 5257
17756 integration 26
17757 integrationen 20
17758 integrationens 2
17759 integrationsfaktor 1
17760 integrationsförfarande 1
17761 integrationsförmåga 1
17762 integrationsmekanismer 1
17763 integrationsmodellen 1
17764 integrationspolitik 3
17765 integrationsproblem 1
17766 integrationsprocess 2
17767 integrationsprocessen 5
17768 integrationsprogram 1
17769 integrationsstrategi 1
17770 integrationsåtgärderna 1
17771 integrera 19
17772 integrerad 15
17773 integrerade 4
17774 integrerades 1
17775 integrerandet 1
17776 integrerar 3
17777 integreras 13
17778 integrerat 5
17779 integrerats 1
17780 integrering 28
17781 integreringen 7
17782 integreringsarbetet 1
17783 integreringsprocesser 1
17784 integritet 6
17785 integriteten 1
17786 intellektuell 3
17787 intellektuella 7
17788 intellektuellt 3
17789 intelligens 2
17790 intelligensen 1
17791 intelligent 8
17792 intelligenta 5
17793 intensifiera 5
17794 intensifieras 1
17795 intensifieringen 1
17796 intensitet 3
17797 intensiteten 1
17798 intensiv 6
17799 intensiva 5
17800 intensivare 1
17801 intensivt 14
17802 intentioner 4
17803 intentionerna 1
17804 inter-etniska 3
17805 interaktiv 3
17806 interaktivitet 2
17807 interaktivitetsnivå 1
17808 interetniska 1
17809 interim 1
17810 interimsavtalen 1
17811 interimsavtalet 4
17812 interimsbetalningar 2
17813 interimsparlament 1
17814 interimspresident 1
17815 interimsråd 2
17816 interimstrukturer 1
17817 interimsåtgärder 1
17818 interinstitutionell 3
17819 interinstitutionella 9
17820 interinstitutionellt 6
17821 intern 14
17822 interna 30
17823 international-socialistiskt 1
17824 internationalisering 1
17825 internationaliseringen 1
17826 internationalistiska 2
17827 internationell 59
17828 internationella 148
17829 internationellt 31
17830 internering 1
17831 interneringar 1
17832 interneringscentra 1
17833 interneringslägret 1
17834 internt 10
17835 interparlamentariska 1
17836 interregionala 4
17837 interregionalt 3
17838 intervall 2
17839 intervaller 3
17840 intervallet 2
17841 intervenera 2
17842 intervenerar 1
17843 intervention 8
17844 interventioner 5
17845 interventionism 2
17846 interventionskapaciteten 1
17847 interventionsrätt 1
17848 interventionsstödet 1
17849 intervju 2
17850 intervjuades 1
17851 intet 8
17852 intetsägande 1
17853 intill 7
17854 intilliggande 2
17855 intima 1
17856 intimt 4
17857 intog 6
17858 intogs 2
17859 intolerans 5
17860 intoleransen 2
17861 intoleransens 2
17862 intolerant 1
17863 intoleranta 2
17864 intonation 1
17865 intranät 2
17866 intressant 36
17867 intressanta 17
17868 intresse 85
17869 intresseföreningar 1
17870 intresseföreningarna 1
17871 intressekonflikter 2
17872 intressemotsättningar 1
17873 intressen 111
17874 intressena 14
17875 intressenter 1
17876 intressera 4
17877 intresserad 13
17878 intresserade 16
17879 intresserar 10
17880 intresserat 2
17881 intresseregister 1
17882 intresseregistret 2
17883 intressesfärer 1
17884 intresset 10
17885 intrigera 1
17886 intrigerade 1
17887 introducera 1
17888 introducerade 1
17889 introducerades 1
17890 introducerar 1
17891 introduceras 2
17892 introducerat 1
17893 introducerats 2
17894 introduktionskursen 1
17895 introduktionskurser 2
17896 introduktionskurserna 1
17897 intryck 21
17898 intrycket 23
17899 inträdde 1
17900 inträde 5
17901 inträdesbiljett 1
17902 inträffa 17
17903 inträffad 1
17904 inträffade 14
17905 inträffar 15
17906 inträffat 18
17907 inträngda 1
17908 intränglingar 1
17909 inträngning 1
17910 inträtt 1
17911 intrång 3
17912 intrånget 1
17913 intyg 1
17914 intyga 3
17915 intäkter 11
17916 intäkterna 2
17917 intäktsanalys 1
17918 intäktsbaserade 1
17919 intäktsförluster 1
17920 intåg 1
17921 inuti 2
17922 invaggade 1
17923 invald 1
17924 invalidiserad 1
17925 invandrad 1
17926 invandrade 7
17927 invandrarbefolkningen 1
17928 invandrare 25
17929 invandrares 1
17930 invandrarförläggningar 1
17931 invandrargrupperna 1
17932 invandrarna 6
17933 invandrarnas 2
17934 invandrarpolitik 1
17935 invandring 16
17936 invandringen 8
17937 invandrings- 1
17938 invandringsfientlig 1
17939 invandringsfrågan 1
17940 invandringsfrågorna 1
17941 invandringspolitik 7
17942 invandringspolitiken 2
17943 invandringspolitikens 1
17944 invandringsrättigheterna 1
17945 invandringstryck 1
17946 invasion 1
17947 invecklad 2
17948 invecklade 4
17949 invecklar 1
17950 invecklat 2
17951 inventarium 1
17952 inventering 1
17953 inverka 2
17954 inverkan 16
17955 inverkar 5
17956 investera 15
17957 investerade 2
17958 investerar 5
17959 investerare 10
17960 investeraren 1
17961 investerarens 1
17962 investerarna 8
17963 investerarnas 2
17964 investerarskydd 1
17965 investeras 2
17966 investerat 1
17967 investerats 1
17968 investering 7
17969 investeringar 65
17970 investeringarna 14
17971 investeringen 3
17972 investeringsbanken 1
17973 investeringsfonden 1
17974 investeringsfonder 2
17975 investeringsfonderna 1
17976 investeringsfondernas 1
17977 investeringsformer 1
17978 investeringsförmågan 1
17979 investeringskapital 1
17980 investeringskostnader 1
17981 investeringskostnaderna 1
17982 investeringsmöjligheterna 2
17983 investeringsnivån 1
17984 investeringsorgan 1
17985 investeringspolitik 1
17986 investeringspolitiken 1
17987 investeringsslag 1
17988 investeringsspektrumet 1
17989 investeringssyfte 1
17990 investeringsteknikernas 1
17991 investeringstjänstedirektivet 1
17992 investeringstjänster 3
17993 investeringsutgifterna 1
17994 investeringsändamål 2
17995 invid 1
17996 inviga 2
17997 invigd 1
17998 invigdes 2
17999 invigning 2
18000 invigningen 2
18001 invigningsceremonin 1
18002 invigningsfesten 1
18003 invirad 1
18004 invit 1
18005 inviterade 2
18006 involvera 2
18007 involverad 1
18008 involverade 10
18009 involverar 1
18010 involveras 3
18011 invända 2
18012 invändning 5
18013 invändningar 17
18014 invändningen 2
18015 invänta 3
18016 inväntar 1
18017 invånare 21
18018 invånarna 13
18019 invånarnas 1
18020 inälvor 2
18021 inåt 4
18022 inövade 1
18023 iordningställande 1
18024 irakisk 1
18025 irakiska 5
18026 iranske 1
18027 irländare 1
18028 irländarna 1
18029 irländsk 7
18030 irländska 17
18031 irländskt 3
18032 ironi 2
18033 ironisera 1
18034 ironisk 1
18035 ironiska 1
18036 ironiskt 3
18037 irra 1
18038 irrationella 1
18039 irrationellt 1
18040 irreducitly 1
18041 irreparabla 2
18042 irrgångar 1
18043 irritation 4
18044 irritationsmoment 1
18045 irriterad 5
18046 irriterade 1
18047 irriterades 1
18048 irriterar 1
18049 irriterat 1
18050 is 4
18051 iscensatt 1
18052 iscensatte 1
18053 isiga 1
18054 iskalla 1
18055 iskallt 1
18056 isolationism 1
18057 isolera 10
18058 isolerad 1
18059 isolerade 6
18060 isoleras 1
18061 isolerat 4
18062 isolering 7
18063 isoleringseffekter 1
18064 israeler 7
18065 israelerna 7
18066 israelisk 2
18067 israelisk-palestinska 1
18068 israeliska 30
18069 israeliske 1
18070 israeliskt 2
18071 issued 3
18072 istapparna 1
18073 istället 6
18074 isvindar 1
18075 isär 7
18076 it 1
18077 italienarna 2
18078 italiensk 4
18079 italienska 34
18080 italienske 2
18081 italienskt 3
18082 iterationer 1
18083 itu 70
18084 iudice 1
18085 iver 4
18086 ivrig 3
18087 ivriga 1
18088 ivrigt 2
18089 iväg 17
18090 iögonenfallande 2
18091 ja 47
18092 jacka 1
18093 jackärmen 1
18094 jag 3499
18095 jagar 3
18096 jakt 8
18097 jakten 3
18098 jaktområdet 1
18099 jakträtt 1
18100 jamaicanska 1
18101 janela 1
18102 januari 60
18103 januarisessionen 1
18104 janushuvud 1
18105 japaner 1
18106 japanska 1
18107 japanskt 1
18108 jargong 2
18109 jargongen 2
18110 jaså 2
18111 jettons 1
18112 jiddisch 5
18113 jingel 1
18114 jingle-belling 1
18115 jobb 39
18116 jobb-med-framtidsutsikter 1
18117 jobba 4
18118 jobbar 3
18119 jobbat 1
18120 jobben 2
18121 jobbet 5
18122 jobbig 1
18123 joint 1
18124 jojo 1
18125 jojoar 1
18126 jojon 3
18127 jokertecken 5
18128 jokertecknen 2
18129 jokertecknet 1
18130 joniserande 1
18131 jord 15
18132 jordaniska 1
18133 jordbruk 35
18134 jordbrukare 17
18135 jordbrukaren 2
18136 jordbrukares 1
18137 jordbrukarfientliga 1
18138 jordbrukarna 7
18139 jordbrukarnas 3
18140 jordbrukarorganisationer 1
18141 jordbruken 3
18142 jordbruket 36
18143 jordbrukets 7
18144 jordbruks 1
18145 jordbruks- 3
18146 jordbruksaktiviteterna 1
18147 jordbruksavsnittet 1
18148 jordbruksbakgrund 1
18149 jordbruksbefolkningen 1
18150 jordbruksekonomin 1
18151 jordbruksexporten 1
18152 jordbruksfonden 1
18153 jordbruksfrågornas 1
18154 jordbruksinkomsterna 2
18155 jordbrukskooperativa 1
18156 jordbrukslobbyn 1
18157 jordbruksmarken 1
18158 jordbruksministern 1
18159 jordbruksmodellen 1
18160 jordbruksnäring 1
18161 jordbruksnäringen 2
18162 jordbruksområden 1
18163 jordbruksområdena 2
18164 jordbruksområdenas 1
18165 jordbruksområdet 2
18166 jordbrukspolitik 9
18167 jordbrukspolitiken 25
18168 jordbrukspraxis 1
18169 jordbrukspriserna 1
18170 jordbruksprodukt 1
18171 jordbruksprodukter 5
18172 jordbruksproduktionen 2
18173 jordbruksreformer 1
18174 jordbruksregionerna 1
18175 jordbrukssektorer 1
18176 jordbrukssektorn 12
18177 jordbrukssektorns 1
18178 jordbrukssynpunkt 1
18179 jordbruksutgifterna 1
18180 jordbruksutskott 1
18181 jordbruksutskottet 1
18182 jordbruksutställningar 1
18183 jordbruksverksamhet 1
18184 jordbävningar 1
18185 jordbävningarna 3
18186 jordbävningen 1
18187 jordbävningsdrabbade 1
18188 jordbävningsdramat 1
18189 jordbävningsfara 2
18190 jordbävningssäkra 1
18191 jordbävningsutsatta 1
18192 jorden 11
18193 jordens 8
18194 jordetunnan 1
18195 jordgubbar 1
18196 jordgubbs- 1
18197 jordiskt 1
18198 jordklotet 1
18199 jordklotets 1
18200 jordluktande 1
18201 jordmån 1
18202 jordnära 1
18203 jordnötsformad 1
18204 jordnötssmörglassar 1
18205 jordskalv 1
18206 jordägare 1
18207 journalismen 1
18208 journalist 2
18209 journalisten 10
18210 journalister 8
18211 journalisterna 5
18212 journalisters 1
18213 journalistiska 1
18214 journalists 2
18215 jovialitet 1
18216 ju 229
18217 jubel 2
18218 jubileumsåret 1
18219 jubla 1
18220 jublande 1
18221 judar 7
18222 judarna 5
18223 judarnas 1
18224 judars 2
18225 jude 7
18226 judegrabbens 1
18227 judeutrotning 1
18228 judisk 3
18229 judiska 7
18230 jugoslaviska 19
18231 jul 3
18232 julen 3
18233 julferien 1
18234 juli 24
18235 julklappar 1
18236 julklappsstämning 1
18237 jultomten 1
18238 jumprar 1
18239 jungfrutal 3
18240 juni 40
18241 jure 2
18242 juridisk 14
18243 juridiska 28
18244 juridiskt 16
18245 juris 7
18246 jurisdiktion 7
18247 jurist 1
18248 jurister 3
18249 juristerna 2
18250 juristlingvisterna 1
18251 just 287
18252 justera 3
18253 justerade 1
18254 justerades 6
18255 justerar 2
18256 justeras 3
18257 justering 1
18258 justeringar 4
18259 justeringsfaktor 1
18260 justice 4
18261 justitie- 1
18262 justitiedepartementet 2
18263 justitieminister 1
18264 justitieministern 1
18265 justitieministerns 1
18266 juveler 1
18267 jäkla 2
18268 jämför 6
18269 jämföra 4
18270 jämförande 1
18271 jämföras 2
18272 jämförbar 1
18273 jämförbara 11
18274 jämförbarhet 1
18275 jämförda 1
18276 jämförelse 13
18277 jämförelsen 1
18278 jämförelser 1
18279 jämförelsevis 1
18280 jämförliga 1
18281 jämförligt 1
18282 jämfört 30
18283 jämka 1
18284 jämlik 2
18285 jämlika 2
18286 jämlikar 1
18287 jämlikhet 15
18288 jämlikheten 6
18289 jämlikhetsperspektiv 1
18290 jämlikt 3
18291 jämmer 1
18292 jämn 6
18293 jämna 3
18294 jämnade 2
18295 jämnan 1
18296 jämnt 3
18297 jämnvikten 1
18298 jämsides 2
18299 jämställande 1
18300 jämställd 3
18301 jämställda 2
18302 jämställde 1
18303 jämställdes 1
18304 jämställdhet 28
18305 jämställdheten 8
18306 jämställdhets- 1
18307 jämställdhetsaspekten 2
18308 jämställdhetsdirektiven 1
18309 jämställdhetsfrågor 10
18310 jämställdhetsfrågorna 1
18311 jämställdhetsperspektiv 2
18312 jämställdhetsperspektivet 1
18313 jämställdhetsplanet 1
18314 jämställdhetstänkande 2
18315 jämställdhetstänkandet 1
18316 jämställdhetsutbildning 2
18317 jämställt 1
18318 jämt 4
18319 jämte 2
18320 jämvikt 10
18321 jämvikten 3
18322 järn- 2
18323 järnindustrin 1
18324 järnkrage 1
18325 järnlängd 1
18326 järnring 1
18327 järnrör 1
18328 järnväg 14
18329 järnvägar 2
18330 järnvägarna 2
18331 järnvägen 6
18332 järnvägens 1
18333 järnvägsföretag 1
18334 järnvägsföretagen 1
18335 järnvägslinjerna 1
18336 järnvägsnät 2
18337 järnvägsnäten 1
18338 järnvägsområde 1
18339 järnvägssektorn 1
18340 järnvägsspår 1
18341 järnvägsövergången 1
18342 järtecken 1
18343 jätte 1
18344 jätteglad 1
18345 jättehårt 1
18346 jättelik 1
18347 jättelikt 1
18348 jätteorder 1
18349 jättestadens 1
18350 jättestor 1
18351 jättestora 2
18352 jättestort 1
18353 jättetankerna 1
18354 jävla 1
18355 k 1
18356 kabarébetonat 1
18357 kabeln 1
18358 kabinen 1
18359 kabinett 2
18360 kabinettet 1
18361 kabinettspost 1
18362 kablar 1
18363 kadaver 1
18364 kadmium 4
18365 kadrer 1
18366 kaffe 4
18367 kaffet 2
18368 kafé 2
18369 kajen 1
18370 kaka 2
18371 kakao 1
18372 kakao- 1
18373 kakaoodlarnas 1
18374 kal 1
18375 kala 1
18376 kalender 1
18377 kalipers 1
18378 kalkrester 1
18379 kalkylblad 2
18380 kalkylbladsliknande 1
18381 kalkyleras 1
18382 kall 2
18383 kalla 43
18384 kallad 12
18385 kallade 47
18386 kallades 5
18387 kallar 19
18388 kallare 1
18389 kallas 15
18390 kallat 13
18391 kallblodiga 1
18392 kallbrun 1
18393 kallelse 1
18394 kallelsen 1
18395 kallsvettig 1
18396 kallt 3
18397 kallvattenarter 1
18398 kalven 1
18399 kam 2
18400 kambodjanska 1
18401 kamera 1
18402 kamma 1
18403 kammar 1
18404 kammare 78
18405 kammaren 91
18406 kammarens 9
18407 kammares 4
18408 kamp 29
18409 kampanj 6
18410 kampanjen 3
18411 kampanjer 2
18412 kampen 45
18413 kamrat 2
18414 kamrater 1
18415 kan 2425
18416 kanadensare 1
18417 kanadensisk 1
18418 kanadensiska 3
18419 kanadensiskt 1
18420 kanal 9
18421 kanalen 2
18422 kanaler 6
18423 kanalerna 1
18424 kanderade 1
18425 kandidat 1
18426 kandidater 5
18427 kandidaterna 3
18428 kandidatland 6
18429 kandidatlandstatus 1
18430 kandidatlista 1
18431 kandidatländer 14
18432 kandidatländerna 25
18433 kandidatländernas 8
18434 kandidatprojekten 1
18435 kandidatur 1
18436 kandiderar 2
18437 kanhända 3
18438 kaninen 1
18439 kaniner 1
18440 kaninunge 1
18441 kanoner 2
18442 kanske 209
18443 kansler 2
18444 kanslern 3
18445 kansli 2
18446 kanslichefer 1
18447 kanslierna 1
18448 kanslisekreteraren 1
18449 kant 2
18450 kanten 3
18451 kanter 1
18452 kantonernas 1
18453 kantstött 1
18454 kaos 6
18455 kaoset 1
18456 kaotisk 1
18457 kapabel 3
18458 kapacitet 25
18459 kapaciteten 4
18460 kapacitetsbyggnad 1
18461 kapacitetsstöd 1
18462 kapacitetsutveckling 1
18463 kapade 1
18464 kapar 1
18465 kapital 17
18466 kapitalbeskattningen 1
18467 kapitalbildning 1
18468 kapitalet 11
18469 kapitalinkomster 4
18470 kapitalinvesteringstillväxt 1
18471 kapitaliseringsförmåga 1
18472 kapitalistiska 4
18473 kapitalkrav 2
18474 kapitalmarknader 1
18475 kapitalmarknaderna 5
18476 kapitalplaceringar 1
18477 kapitalrörelser 1
18478 kapitalskatt 3
18479 kapitalskatter 1
18480 kapitaltillskott 1
18481 kapitalutnyttjande 1
18482 kapitel 19
18483 kapitelrubrikerna 1
18484 kapitlet 3
18485 kapitulera 1
18486 kapitulerar 1
18487 kapp 2
18488 kapplöpningshaj 1
18489 kapsyler 1
18490 kapten 3
18491 kaptenen 2
18492 kaptener 1
18493 karaff 1
18494 karakteriserade 1
18495 karakteriserar 1
18496 karakteriseringar 1
18497 karakteristisk 1
18498 karakteristiska 1
18499 karakteristiskt 3
18500 karaktär 32
18501 karaktären 8
18502 karaktärer 1
18503 karaktäristisk 1
18504 kareernas 1
18505 karga 2
18506 karikatyr 1
18507 karl 3
18508 karlar 1
18509 karmosinröd 1
18510 karriärer 1
18511 karriärmöjligheter 1
18512 karriärplanering 1
18513 karriärstegen 1
18514 karta 1
18515 kartan 5
18516 kartell- 3
18517 kartellbestämmelserna 1
18518 kartellbildningar 1
18519 karteller 1
18520 kartellförbudet 2
18521 kartellmyndighet 1
18522 kartellrätten 4
18523 kartlägger 1
18524 kartläggning 3
18525 kartonger 1
18526 kartor 3
18527 kasino 2
18528 kaskad 1
18529 kassa 1
18530 kassaapparaten 1
18531 kasserade 3
18532 kassettband 1
18533 kasta 4
18534 kastade 10
18535 kastades 3
18536 kastar 3
18537 kastas 4
18538 kastat 1
18539 kastats 1
18540 kastvapen 1
18541 katalog 4
18542 katalogens 1
18543 katalysator 3
18544 katalytisk 1
18545 katastrof 43
18546 katastrofala 8
18547 katastrofberedskap 1
18548 katastrofdrabbade 3
18549 katastrofen 29
18550 katastrofens 2
18551 katastrofer 34
18552 katastroferna 5
18553 katastrofhjälp 2
18554 katastrofplatsen 1
18555 katastrofprogram 1
18556 katastrofsituation 1
18557 katastrofsituationen 1
18558 katastrofstrategi 1
18559 katastrofstöd 2
18560 kategori 5
18561 kategorier 7
18562 kategorierna 4
18563 kategorifält 3
18564 kategorifältområde 1
18565 kategoriska 1
18566 kategoriskt 1
18567 katolicismen 1
18568 katolik 2
18569 katoliker 3
18570 katolikernas 1
18571 katolska 5
18572 katt 1
18573 katter 1
18574 kattflatan 1
18575 kattlapp 1
18576 kattliknande 1
18577 kattun 1
18578 kattuntryck 1
18579 kavaj 1
18580 kavaljerer 1
18581 kedja 5
18582 kedjan 5
18583 kedjefångarna 1
18584 kedjorna 1
18585 kejsardömets 1
18586 kejsaren 1
18587 keltiska 2
18588 kemiindustrins 1
18589 kemikalier 9
18590 kemikaliestrategin 1
18591 kemisk 2
18592 kemiska 13
18593 kerubliknande 1
18594 kex 1
18595 kg 2
18596 khakishorts 1
18597 khmererna 2
18598 khmerernas 2
18599 kibbutzen 2
18600 kibbutzsjöman 1
18601 kick 1
18602 kidnappningar 1
18603 kika 1
18604 kikade 1
18605 kil 1
18606 kila 1
18607 kilar 1
18608 kilo 5
18609 kilometer 8
18610 kilowattimme 1
18611 kind 1
18612 kinden 1
18613 kinder 2
18614 kinderna 1
18615 kindknotor 1
18616 kineser 1
18617 kineserna 3
18618 kinesisk 1
18619 kinesiska 18
18620 kinesiskt 1
18621 kinkig 1
18622 kirurgiskt 1
18623 kisade 1
18624 kista 1
18625 kittel 1
18626 kitteln 1
18627 kjolarna 1
18628 kl 1
18629 kl. 92
18630 kl.12.00 1
18631 klackar 1
18632 kladdade 1
18633 klaga 1
18634 klagade 1
18635 klagan 1
18636 klagar 2
18637 klagat 1
18638 klagoandar 1
18639 klagomål 15
18640 klagomålet 2
18641 klagomålsförfarande 1
18642 klagoskrivelse 1
18643 klagosånger 1
18644 klamrande 2
18645 klandervärt 1
18646 klandras 2
18647 klanen 1
18648 klappa 1
18649 klappade 1
18650 klappjakt 1
18651 klar 44
18652 klara 54
18653 klarade 4
18654 klarades 1
18655 klarar 17
18656 klarare 2
18657 klaras 1
18658 klarast 1
18659 klarat 2
18660 klarats 1
18661 klargjorde 1
18662 klargjordes 1
18663 klargjort 8
18664 klargör 10
18665 klargöra 25
18666 klargörande 7
18667 klargöranden 3
18668 klargörandet 1
18669 klargöras 4
18670 klargörs 8
18671 klarhet 15
18672 klarheten 1
18673 klarhetens 1
18674 klarlagd 1
18675 klarlagt 1
18676 klarlagts 1
18677 klarlägga 3
18678 klarläggande 4
18679 klarlägganden 2
18680 klarläggandena 1
18681 klarläggandet 1
18682 klarläggas 1
18683 klarsynthet 1
18684 klart 168
18685 klartecken 5
18686 klartext 7
18687 klass 6
18688 klassa 1
18689 klassas 1
18690 klassats 1
18691 klassen 3
18692 klassens 1
18693 klasser 1
18694 klassernas 1
18695 klassificera 3
18696 klassificerar 1
18697 klassificerat 2
18698 klassificering 1
18699 klassificeringen 1
18700 klassificeringsbolagen 1
18701 klassificeringsregister 1
18702 klassificeringssällskapen 4
18703 klassificeringssällskapet 1
18704 klassisk 1
18705 klassiska 5
18706 klassiskt 3
18707 klausul 4
18708 klausulen 2
18709 klausuler 5
18710 klaveret 1
18711 klen 1
18712 klent 1
18713 klev 8
18714 kliande 1
18715 klibbiga 2
18716 klick 2
18717 klient 1
18718 klienter 2
18719 klientilism 1
18720 klimat 13
18721 klimatet 11
18722 klimatfrågor 1
18723 klimatförändring 2
18724 klimatförändringar 5
18725 klimatförändringarna 3
18726 klimatförändringen 2
18727 klimatiska 2
18728 klimatmässiga 1
18729 klimatmönster 1
18730 klimatologiska 2
18731 klimatprotokoll 1
18732 klimatskillnader 1
18733 klingande 2
18734 kliniska 1
18735 kliniskt 1
18736 klippan 1
18737 klippas 1
18738 klippblock 2
18739 klippbranten 1
18740 klippkaos 1
18741 klippstup 1
18742 klippte 2
18743 klirr 1
18744 klirret 1
18745 klistra 1
18746 klistrat 1
18747 kliv 2
18748 kliver 1
18749 kloaklukt 1
18750 klocka 1
18751 klocka-bracelet 1
18752 klockan 15
18753 klok 7
18754 kloka 2
18755 klokare 2
18756 klokast 1
18757 klokhet 1
18758 klokt 20
18759 klon 1
18760 klorna 1
18761 kloten 1
18762 klotter 1
18763 klumparna 1
18764 klungor 2
18765 klunk 1
18766 klunkar 1
18767 kluven 1
18768 kluvenhet 1
18769 klyfta 2
18770 klyftan 7
18771 klyftor 2
18772 klyftorna 3
18773 klyva 1
18774 klä 2
18775 kläckts 1
18776 klädborste 1
18777 klädd 5
18778 klädda 2
18779 klädde 1
18780 kläder 14
18781 kläderna 2
18782 klädnad 1
18783 klädnader 2
18784 klämde 3
18785 klänning 4
18786 klätt 1
18787 klättra 2
18788 klättrade 4
18789 km 5
18790 knacka 1
18791 knackade 1
18792 knackat 1
18793 knall 1
18794 knallrött 1
18795 knapp 5
18796 knappa 5
18797 knappar 1
18798 knappast 31
18799 knappen 2
18800 knappnålshuvuden 1
18801 knappt 16
18802 knarrar 1
18803 knaster 1
18804 knastrade 1
18805 knep 2
18806 knepiga 1
18807 knipa 1
18808 kniv 2
18809 knivar 2
18810 knivarnas 1
18811 knivhuggen 2
18812 knogande 1
18813 knollrigt 1
18814 knoppigt 1
18815 knorvig 1
18816 knotande 1
18817 know-how 3
18818 knubbig 1
18819 knuff 1
18820 knuffa 1
18821 knuffade 2
18822 knussla 1
18823 knuten 6
18824 knutet 3
18825 knutna 9
18826 knutpunkt 1
18827 knutpunkterna 1
18828 knyckte 1
18829 knyta 10
18830 knytas 2
18831 knyter 3
18832 knyts 1
18833 knä 4
18834 knäcka 1
18835 knäckas 1
18836 knäckt 1
18837 knäckte 2
18838 knän 1
18839 knäna 4
18840 knäppklocka 1
18841 knät 1
18842 knåpat 1
18843 knölar 1
18844 knöt 1
18845 ko 2
18846 ko-affären 1
18847 ko-krisen 1
18848 koalition 3
18849 koalitionen 3
18850 koalitionens 2
18851 koalitionsavtalen 1
18852 koalitionsförhandlingarna 2
18853 koalitionsregering 4
18854 koalitionssamtal 1
18855 kock 2
18856 kockmössa 1
18857 kod 2
18858 koden 3
18859 koder 1
18860 kodifiera 1
18861 kodifierad 3
18862 kodifieras 1
18863 kodifikationen 1
18864 koffertar 1
18865 kofferten 4
18866 koherens 1
18867 koherensen 1
18868 kokade 1
18869 kokhett 1
18870 kokong 1
18871 kokor 1
18872 kokosnötterna 1
18873 kol 1
18874 kol- 1
18875 koldioxid 5
18876 koldioxiden 1
18877 koldioxidskatt 1
18878 koldioxidutsläppen 1
18879 koleldad 1
18880 kolera 1
18881 kolförrådet 1
18882 kolhög 1
18883 kolja 2
18884 kollaps 3
18885 kollapsa 2
18886 kollega 124
18887 kollegan 26
18888 kollegans 1
18889 kollegas 3
18890 kolleger 266
18891 kollegerna 21
18892 kollegernas 4
18893 kollegers 8
18894 kollegiala 1
18895 kollegialiteten 1
18896 kollegiet 1
18897 kollegium 2
18898 kollegor 32
18899 kollegorna 1
18900 kollegors 4
18901 kollektiv 3
18902 kollektiva 17
18903 kollektivavtal 7
18904 kollektivet 1
18905 kollektivt 2
18906 kollektivtrafik 1
18907 kollektivtrafiken 1
18908 kollisioner 1
18909 kollisionskurs 2
18910 koloni 1
18911 koloniala 2
18912 kolonialdepartementet 1
18913 kolonialdepartementets 1
18914 kolonialism 1
18915 kolonialister 1
18916 kolonialisterna 1
18917 kolonialmakterna 1
18918 kolonialtiden 1
18919 kolonialtjänsteman 2
18920 kolonialtjänstemännen 1
18921 kolonialtyp 1
18922 kolonier 2
18923 kolonisatörer 3
18924 kolonist 1
18925 kolonisterna 1
18926 koloss 1
18927 kolossala 2
18928 kolossalt 4
18929 kolumn- 2
18930 kolumner 1
18931 kolumnerna 1
18932 kolumnfält 2
18933 kolumnnamn 2
18934 kolumnområden 1
18935 kolumnområdet 1
18936 kolväten 1
18937 kom 158
18938 kombination 9
18939 kombinationen 1
18940 kombinationer 1
18941 kombinera 3
18942 kombinerade 1
18943 kombinerar 3
18944 kombineras 3
18945 kombinerat 1
18946 komedi 1
18947 komet 1
18948 kometen 1
18949 kometerna 1
18950 komisk 1
18951 komissionen 2
18952 komma 280
18953 komma-av-åldern 1
18954 kommande 123
18955 kommandon 1
18956 kommandostyrkor 2
18957 kommandot 8
18958 kommas 1
18959 kommen 1
18960 kommendera 1
18961 kommentar 15
18962 kommentarer 36
18963 kommentarerna 4
18964 kommentarsblock 1
18965 kommentatorers 1
18966 kommentera 22
18967 kommenterades 1
18968 kommenterat 1
18969 kommer 1957
18970 kommers 1
18971 kommersiell 5
18972 kommersiella 14
18973 kommersiellt 4
18974 kommission 48
18975 kommissionen 1437
18976 kommissionens 463
18977 kommissionsakt 1
18978 kommissionsdirektoratet 1
18979 kommissionsförslag 1
18980 kommissionskollegiet 1
18981 kommissionsledamot 6
18982 kommissionsledamoten 8
18983 kommissionsledamöter 4
18984 kommissionsledamöterna 3
18985 kommissionsledamöters 1
18986 kommissionsnivå 1
18987 kommissionsordförande 34
18988 kommissionsordföranden 1
18989 kommissionssystemet 1
18990 kommissionstjänsten 1
18991 kommissionär 457
18992 kommissionären 120
18993 kommissionärens 9
18994 kommissionärer 28
18995 kommissionärerna 13
18996 kommissionärernas 2
18997 kommissionärs 1
18998 kommissionärskolleger 1
18999 kommit 100
19000 kommitté 12
19001 kommittédjungel 1
19002 kommittéer 7
19003 kommittéerna 8
19004 kommittéförfarande 2
19005 kommittéförfaranden 6
19006 kommittéförfarandena 2
19007 kommittéförfarandesystemet 2
19008 kommittéförfarandet 16
19009 kommittén 15
19010 kommitténs 1
19011 kommittésystemet 2
19012 kommun 2
19013 kommunal 3
19014 kommunala 7
19015 kommunalparlament 1
19016 kommuner 7
19017 kommunerna 4
19018 kommunfullmäktige 3
19019 kommunicera 1
19020 kommunicerande 1
19021 kommunicerar 1
19022 kommunicerat 1
19023 kommunikation 9
19024 kommunikationen 4
19025 kommunikationer 6
19026 kommunikationerna 1
19027 kommunikations- 1
19028 kommunikationskampanj 1
19029 kommunikationskanaler 2
19030 kommunikationsklyftan 1
19031 kommunikationsmedlen 2
19032 kommunikationsområdet 1
19033 kommunikationsproblemet 1
19034 kommunikationsstrategi 1
19035 kommunikationsteknik 1
19036 kommunikationstekniken 1
19037 kommunikationstjänster 1
19038 kommuniké 1
19039 kommunikéer 1
19040 kommunism 2
19041 kommunismen 2
19042 kommunismens 2
19043 kommunisterna 2
19044 kommunistiska 4
19045 kommunistiskt 2
19046 kommunistpartis 1
19047 kommunistregimerna 1
19048 kommunvalen 1
19049 kompakta 1
19050 kompaniets 1
19051 kompass 1
19052 kompatibelt 2
19053 kompatibla 2
19054 kompensation 17
19055 kompensationer 2
19056 kompensationsfonderna 1
19057 kompensationsåtgärden 1
19058 kompensationsåtgärder 2
19059 kompensationsåtgärderna 2
19060 kompensera 7
19061 kompenserade 1
19062 kompenserades 1
19063 kompenserande 1
19064 kompenserar 3
19065 kompenseras 3
19066 kompenserats 1
19067 kompetens 24
19068 kompetensen 3
19069 kompetenskrav 1
19070 kompetensområden 2
19071 kompetent 8
19072 kompetenta 3
19073 kompisar 1
19074 komplement 15
19075 komplementaritet 2
19076 komplementaritetsprinciperna 1
19077 komplett 5
19078 komplettera 23
19079 kompletterad 1
19080 kompletterande 18
19081 kompletterar 5
19082 kompletteras 4
19083 kompletterat 1
19084 komplettering 5
19085 komplex 1
19086 komplexa 5
19087 komplexitet 3
19088 komplexiteten 1
19089 komplext 5
19090 komplicerad 17
19091 komplicerade 12
19092 komplicerar 1
19093 komplicerat 19
19094 komplikationer 3
19095 komplimang 1
19096 komplimanger 10
19097 komplimentera 1
19098 komplotter 1
19099 komponent 2
19100 komponenten 1
19101 komponenter 8
19102 komponenterna 15
19103 komposteringen 1
19104 kompromettera 1
19105 kompromiss 24
19106 kompromissa 5
19107 kompromissa.§ 1
19108 kompromissarbete 1
19109 kompromissen 5
19110 kompromisser 6
19111 kompromissförslag 4
19112 kompromisslös 1
19113 kompromisslöshet 1
19114 kompromisslösheten 2
19115 kompromisslösning 5
19116 kompromissresolution 1
19117 kompromissresolutionen 4
19118 kompromissrundan 1
19119 kompromisstexten 1
19120 koncentration 14
19121 koncentrationen 6
19122 koncentrationer 7
19123 koncentrationsläger 2
19124 koncentrationslägren 1
19125 koncentrationslägrens 1
19126 koncentrationsprincipen 1
19127 koncentrera 34
19128 koncentrerad 3
19129 koncentrerade 1
19130 koncentrerar 10
19131 koncentreras 7
19132 koncentrerat 5
19133 koncentrerats 1
19134 koncentrisk 1
19135 koncept 10
19136 konceptet 5
19137 koncern 1
19138 koncerner 1
19139 koncis 2
19140 koncisa 1
19141 koncist 2
19142 kondition 1
19143 konfederal 1
19144 konfederation 1
19145 konferens 15
19146 konferensen 21
19147 konferensens 1
19148 konferenserna 3
19149 konfession 1
19150 konfessionslöst 1
19151 konfidentiell 1
19152 konfidentiella 3
19153 konfigurerar 1
19154 konfiskera 1
19155 konfiskerad 1
19156 konfiskerats 1
19157 konflikt 18
19158 konflikten 19
19159 konfliktens 1
19160 konflikter 34
19161 konflikterna 3
19162 konfliktförebyggande 13
19163 konflikthantering 2
19164 konfliktlösning 7
19165 konfliktorsakande 1
19166 konformism 1
19167 konfrontation 1
19168 konfrontationer 1
19169 konfrontationspolitik 1
19170 konfrontera 1
19171 konfronterades 1
19172 konfronteras 7
19173 kongolesisk 1
19174 kongolesiska 1
19175 kongotyg 1
19176 kongress 1
19177 kongressen 2
19178 kongressmän 1
19179 konjaksglasen 1
19180 konjaksglaset 1
19181 konjunktur 1
19182 konjunkturberoende 1
19183 konjunkturbetingad 1
19184 konjunkturcykeln 1
19185 konjunkturen 3
19186 konjunkturer 1
19187 konjunkturmässiga 1
19188 konjunkturmässigt 1
19189 konjunktursituation 1
19190 konjunktursvängningarna 1
19191 konkret 63
19192 konkreta 104
19193 konkretare 1
19194 konkretaste 1
19195 konkretisera 7
19196 konkretiserar 1
19197 konkretiseras 3
19198 konkretiserats 1
19199 konkretisering 1
19200 konkretiseringar 1
19201 konkurrens 83
19202 konkurrens- 2
19203 konkurrensaspekten 1
19204 konkurrensavgöranden 1
19205 konkurrensbegränsande 2
19206 konkurrensbegränsningar 1
19207 konkurrensbestämmelser 4
19208 konkurrensbestämmelserna 2
19209 konkurrensdebatt 1
19210 konkurrensdebatten 1
19211 konkurrensdomstol 1
19212 konkurrensdugliga 1
19213 konkurrensduglighet 1
19214 konkurrensen 80
19215 konkurrensens 3
19216 konkurrensfriheten 1
19217 konkurrensfrämjande 1
19218 konkurrensfråga 1
19219 konkurrensfrågan 1
19220 konkurrensfrågor 2
19221 konkurrensfrågorna 2
19222 konkurrensfördel 2
19223 konkurrensfördelar 1
19224 konkurrensförfarandet 1
19225 konkurrensförmåga 2
19226 konkurrensförmågan 1
19227 konkurrenshinder 2
19228 konkurrenshämmande 2
19229 konkurrensinitiativen 1
19230 konkurrensinriktad 1
19231 konkurrensjämvikt 1
19232 konkurrenskraft 34
19233 konkurrenskraften 18
19234 konkurrenskraftens 1
19235 konkurrenskraftig 11
19236 konkurrenskraftiga 16
19237 konkurrenskraftigare 2
19238 konkurrenskraftigaste 1
19239 konkurrenskraftigt 2
19240 konkurrenskriterier 1
19241 konkurrenskriterierna 1
19242 konkurrenskultur 3
19243 konkurrenskulturens 1
19244 konkurrenskulturerna 1
19245 konkurrensmedel 1
19246 konkurrensminister 1
19247 konkurrensmyndighet 3
19248 konkurrensmyndigheten 1
19249 konkurrensmyndigheterna 3
19250 konkurrensmyndigheternas 1
19251 konkurrensmyndigheters 1
19252 konkurrensmål 1
19253 konkurrensmöjligheter 1
19254 konkurrensnackdel 1
19255 konkurrensnackdelen 1
19256 konkurrensområdet 3
19257 konkurrensordning 1
19258 konkurrenspakter 1
19259 konkurrenspolitik 20
19260 konkurrenspolitiken 41
19261 konkurrenspolitikens 6
19262 konkurrenspolitisk 1
19263 konkurrenspolitiska 3
19264 konkurrenspolitiskt 2
19265 konkurrensprincipen 3
19266 konkurrenspräglad 1
19267 konkurrensregler 1
19268 konkurrensreglerna 9
19269 konkurrensrelaterade 1
19270 konkurrensrätt 1
19271 konkurrensrätten 6
19272 konkurrensrättens 1
19273 konkurrensrättsliga 1
19274 konkurrenssituationer 1
19275 konkurrensskadlig 1
19276 konkurrensskyddet 2
19277 konkurrensskäl 1
19278 konkurrensstrid 1
19279 konkurrensstörningar 2
19280 konkurrenssvårigheter 1
19281 konkurrenssynpunkt 1
19282 konkurrenstrycket 1
19283 konkurrensutsatt 1
19284 konkurrensutsätta 2
19285 konkurrensutsättning 1
19286 konkurrensutsättningar 1
19287 konkurrensutsättningen 1
19288 konkurrensverken 1
19289 konkurrensvillkor 5
19290 konkurrensvillkoren 7
19291 konkurrensvänligare 1
19292 konkurrensärenden 2
19293 konkurrent 2
19294 konkurrenter 7
19295 konkurrentländer 1
19296 konkurrera 11
19297 konkurrerar 1
19298 konkurs 3
19299 konkurser 5
19300 konkursfond 1
19301 konsekvens 16
19302 konsekvensen 3
19303 konsekvenser 64
19304 konsekvenserna 36
19305 konsekvensutredning 2
19306 konsekvensutredningar 2
19307 konsekvensutredningarnas 1
19308 konsekvent 28
19309 konsekventa 9
19310 konsensus 2
19311 konsert 1
19312 konserten 1
19313 konservativa 13
19314 konservativas 1
19315 konserver 1
19316 konsolidera 1
19317 konsoliderade 1
19318 konsoliderar 1
19319 konsoliderat 1
19320 konsolidering 5
19321 konsolideringen 3
19322 konsolideringsprogram 1
19323 konsortierna 1
19324 konsortiet 1
19325 konspirationer 1
19326 konst 5
19327 konstant 4
19328 konstatera 69
19329 konstaterade 5
19330 konstaterades 2
19331 konstaterande 4
19332 konstaterandet 2
19333 konstaterar 13
19334 konstateras 4
19335 konstaterat 7
19336 konstaterats 1
19337 konsten 1
19338 konstfullt 1
19339 konstföremål 1
19340 konstgjord 2
19341 konstgjorda 1
19342 konstgjort 1
19343 konstgrepp 1
19344 konstgödsel 1
19345 konstig 1
19346 konstiga 4
19347 konstigt 7
19348 konstituera 1
19349 konstituerades 1
19350 konstitution 5
19351 konstitutionell 4
19352 konstitutionella 23
19353 konstitutionen 1
19354 konstitutivt 1
19355 konstkommittén 1
19356 konstkritikern 1
19357 konstlade 1
19358 konstlat 1
19359 konstlöst 1
19360 konstmuseum 1
19361 konstnären 1
19362 konstnärer 6
19363 konstnärerna 4
19364 konstnärers 4
19365 konstnärliga 3
19366 konstruera 6
19367 konstruerades 1
19368 konstruerat 1
19369 konstruerats 1
19370 konstruktion 9
19371 konstruktionen 1
19372 konstruktioner 1
19373 konstruktionsarbete 1
19374 konstruktionsarbetet 5
19375 konstruktiv 9
19376 konstruktiva 15
19377 konstruktivt 12
19378 konstruktören 1
19379 konstruktörerna 1
19380 konststycken 1
19381 konstverk 1
19382 konsultationer 3
19383 konsultbasis 1
19384 konsulter 1
19385 konsulterande 1
19386 konsulteras 1
19387 konsument 2
19388 konsumenten 16
19389 konsumenten-medborgaren 1
19390 konsumenter 16
19391 konsumenterna 32
19392 konsumenternas 25
19393 konsumenters 1
19394 konsumentfrågor 20
19395 konsumentförtroende 1
19396 konsumentorganisationen 1
19397 konsumentpolitik 4
19398 konsumentpolitisk 1
19399 konsumentrelaterad 1
19400 konsumenträtten 1
19401 konsumentskydd 11
19402 konsumentskyddet 6
19403 konsumentskyddsorganisationerna 1
19404 konsumenttillvänt 1
19405 konsumentvaror 1
19406 konsumentvänligt 1
19407 konsumeras 1
19408 konsumtion 4
19409 konsumtionen 2
19410 kontakt 20
19411 kontaktade 1
19412 kontaktat 3
19413 kontakten 5
19414 kontakter 23
19415 kontakterna 5
19416 kontamination 1
19417 kontaminerade 1
19418 kontanter 1
19419 kontexten 1
19420 kontinent 9
19421 kontinentala 3
19422 kontinentaleuropéerna 1
19423 kontinentalt 1
19424 kontinenten 7
19425 kontinentens 3
19426 kontinenter 1
19427 kontinenterna 1
19428 kontinents 2
19429 kontinuerlig 3
19430 kontinuerligt 5
19431 kontinuitet 3
19432 kontinuiteten 3
19433 konto 1
19434 kontonamnet 1
19435 kontor 11
19436 kontoren 1
19437 kontoret 2
19438 kontorister 1
19439 kontorslokaler 1
19440 kontrahenterna 1
19441 kontrakt 11
19442 kontraktet 2
19443 kontrakts- 1
19444 kontraktsramar 1
19445 kontraktsåtagande 1
19446 kontraproduktiv 1
19447 kontraproduktivt 3
19448 kontrast 3
19449 kontrasten 1
19450 kontraster 1
19451 kontrasterar 1
19452 kontroll 136
19453 kontroll- 2
19454 kontrollanterna 1
19455 kontrollapparat 1
19456 kontrollen 32
19457 kontroller 52
19458 kontrollera 44
19459 kontrollerad 5
19460 kontrollerade 3
19461 kontrollerades 1
19462 kontrollerar 9
19463 kontrolleras 19
19464 kontrollerat 1
19465 kontrollerbara 1
19466 kontrollerna 9
19467 kontrollfunktion 1
19468 kontrollförfarande 1
19469 kontrollförfaranden 2
19470 kontrollförfarandet 1
19471 kontrollmakt 1
19472 kontrollmakten 1
19473 kontrollmedlen 1
19474 kontrollmekanismer 3
19475 kontrollmyndighet 1
19476 kontrollmyndigheterna 1
19477 kontrollmöjlighet 1
19478 kontrollmöjligheter 3
19479 kontrollnamn 1
19480 kontrollnormerna 1
19481 kontrollområdet 1
19482 kontrollorgan 2
19483 kontrollprocessen 1
19484 kontrollprogram 1
19485 kontrollprogrammen 1
19486 kontrollrättigheter 1
19487 kontrollstyrka 1
19488 kontrollsystem 2
19489 kontrollsystemet 1
19490 kontrollsystemets 1
19491 kontrolluppdrag 1
19492 kontrollverksamheten 1
19493 kontrolläger 1
19494 kontrollåtgärder 2
19495 kontrovers 2
19496 kontroversen 2
19497 kontroverser 3
19498 kontroversiell 4
19499 kontroversiella 2
19500 kontroversiellt 4
19501 konturlösa 1
19502 konungariket 1
19503 konvenansflagg 1
19504 konvent 2
19505 konventet 3
19506 konvention 23
19507 konventionell 1
19508 konventionella 3
19509 konventionen 38
19510 konventionens 2
19511 konventioner 13
19512 konventionerna 1
19513 konventionsinstrumenten 1
19514 konventionsnivå 1
19515 konvergens 20
19516 konvergensen 9
19517 konvergenskriterier 6
19518 konvergenskriterierna 3
19519 konvergenskriterium 2
19520 konvergensperspektiv 1
19521 konvergensprocess 1
19522 konvergensprogrammen 1
19523 konvergensstrategi 1
19524 konvergensstrategier 1
19525 konvergensstrategin 1
19526 konvergering 1
19527 konvergeringsprocess 1
19528 konversation 1
19529 konversationen 1
19530 konverserade 1
19531 konvertera 4
19532 konverterade 2
19533 konverteras 3
19534 kooperationens 1
19535 kooperativ 1
19536 kooperativa 1
19537 kopia 4
19538 kopian 1
19539 kopiera 4
19540 kopierade 3
19541 kopierar 5
19542 kopieras 2
19543 kopiering 4
19544 kopieringsrätten 1
19545 kopieringsskyddet 1
19546 kopior 3
19547 kopp 2
19548 koppar 1
19549 kopparbrunt 1
19550 koppen 2
19551 koppla 4
19552 kopplad 5
19553 kopplas 5
19554 kopplat 3
19555 kopplats 1
19556 koppling 8
19557 kopplingarna 1
19558 kopplingen 4
19559 kor 1
19560 kor. 1
19561 korgar 1
19562 korken 1
19563 korna 1
19564 korporatism 1
19565 korpsvart 1
19566 korpus 1
19567 korrekt 44
19568 korrekta 11
19569 korrektare 2
19570 korrekthet 1
19571 korrespondens 1
19572 korrespondent 1
19573 korrespondenten 1
19574 korrespondenter 1
19575 korridoren 1
19576 korridorer 3
19577 korridorerna 1
19578 korridorernas 1
19579 korrigerande 1
19580 korrigeras 2
19581 korrugerad 1
19582 korrumpera 1
19583 korrumperat 2
19584 korrupt 1
19585 korrupta 1
19586 korruption 14
19587 korruptionen 9
19588 korruptionsaffärer 3
19589 korruptionsdömt 1
19590 korruptionsskandal 1
19591 korruptionsskandalerna 1
19592 kors 2
19593 korsade 3
19594 korsar 1
19595 korseld 1
19596 korselden 1
19597 korset 2
19598 korsett 1
19599 korsfråga 4
19600 korslagda 1
19601 korsriddarna 1
19602 kort 134
19603 korta 19
19604 kortare 6
19605 kortas 3
19606 kortaste 1
19607 korten 2
19608 kortet 7
19609 kortets 3
19610 kortfattad 1
19611 kortfattat 2
19612 korthet 3
19613 kortlek 1
19614 kortlivad 2
19615 kortsiktig 2
19616 kortsiktiga 4
19617 kortsiktighet 2
19618 kortsiktigt 2
19619 kortsnaggade 1
19620 kortvarig 1
19621 kortväxt 2
19622 korvar 1
19623 koscherlunch 2
19624 koschermat 2
19625 koschersmörgåsar 1
19626 kosmetika 1
19627 kosovanska 1
19628 kosovoalbaner 6
19629 kosovoalbanerna 3
19630 kosovoalbanska 2
19631 kosta 4
19632 kostade 5
19633 kostar 14
19634 kostat 3
19635 kosthållning 1
19636 kostnad 14
19637 kostnaden 26
19638 kostnader 59
19639 kostnaderna 61
19640 kostnads 1
19641 kostnads- 1
19642 kostnads-intäktsanalys 1
19643 kostnads-intäktsanalysen 1
19644 kostnads-nytto-analys 1
19645 kostnadsbefrielse 1
19646 kostnadsbefrielsen 3
19647 kostnadseffektiv 2
19648 kostnadseffektiva 2
19649 kostnadseffektivt 1
19650 kostnadselementet 1
19651 kostnadsfri 3
19652 kostnadsfria 1
19653 kostnadsfritt 1
19654 kostnadsfördelningen 1
19655 kostnadsinflation 1
19656 kostnadsintensiv 1
19657 kostnadsintensivt 1
19658 kostnadskontroll 1
19659 kostnadspolicy 1
19660 kostnadssystem 4
19661 kostnadstäckande 1
19662 kostnadstäckning 1
19663 kostnadsuppskattning 1
19664 kostnadsutvecklingen 1
19665 kostsam 1
19666 kostsamma 1
19667 kostsamt 3
19668 kostym 4
19669 kostymen 1
19670 kovändning 1
19671 krafsar 1
19672 kraft 87
19673 kraften 11
19674 krafter 16
19675 krafterna 4
19676 krafters 1
19677 kraftfull 6
19678 kraftfulla 10
19679 kraftfullare 2
19680 kraftfullt 16
19681 kraftig 15
19682 kraftiga 8
19683 kraftigare 4
19684 kraftigaste 1
19685 kraftigt 31
19686 kraftmätning 1
19687 kraftnät 1
19688 krafttag 3
19689 kraftåtgärder 1
19690 kragar 3
19691 kragar-ben 1
19692 krage 1
19693 kragen 1
19694 kramade 1
19695 kramat 1
19696 krampen 1
19697 kran 1
19698 kranarna 1
19699 kranin 1
19700 krasande 1
19701 krasch 1
19702 kraschade 1
19703 kraschat 1
19704 krasst 1
19705 krav 119
19706 kravallpoliser 1
19707 kravat 1
19708 kraven 37
19709 kravet 31
19710 kravla 1
19711 kreativ 2
19712 kreativa 5
19713 kreativitet 1
19714 kreativiteten 3
19715 kreativt 1
19716 kreatörer 1
19717 krediter 1
19718 krediterna 1
19719 kreditinstitut 1
19720 kreditvärdighet 2
19721 kreditvärdighetsskala 1
19722 kretensare 1
19723 krets 1
19724 kretsar 3
19725 kretsat 1
19726 kretsen 2
19727 kretslopp 3
19728 krig 48
19729 kriga 2
19730 krigare 1
19731 krigat 1
19732 krigen 2
19733 kriget 30
19734 krigföring 2
19735 krigisk 2
19736 krigsekonomi 1
19737 krigsfartyg 1
19738 krigsflyktingar 1
19739 krigsfångar 1
19740 krigsförbrytardomstolen 1
19741 krigsförbrytare 1
19742 krigsförbrytarförbundets 1
19743 krigsförbrytartribunalen 4
19744 krigsförbrytelser 1
19745 krigsförklaring 1
19746 krigshandlingar 1
19747 krigshandlingarna 1
19748 krigsherrarna 1
19749 krigshärjade 1
19750 krigsivrare 1
19751 krigskonstens 1
19752 krigskorrespondenten 1
19753 krigsmaskin 1
19754 krigsmateriel 1
19755 krigsmålad 1
19756 krigspropagandan 1
19757 krigssituationer 1
19758 krigsskador 1
19759 krigsslutet 1
19760 krigsterminalen 1
19761 krigsutbrott 1
19762 krigsåren 1
19763 kriminalisera 2
19764 kriminaliseras 1
19765 kriminalitet 9
19766 kriminalitetsbekämpning 1
19767 kriminalpolitik 1
19768 kriminalvården 1
19769 kriminell 1
19770 kriminella 5
19771 kriminellt 1
19772 kring 51
19773 kringgå 3
19774 kringgående 2
19775 kringgår 1
19776 kringgås 1
19777 kringirrande 1
19778 kringliggande 1
19779 kringskuren 1
19780 kringskuret 1
19781 kringspridda 1
19782 kringströvanden 1
19783 kringvärvd 1
19784 kringvärvde 1
19785 kris 19
19786 krisbildningarna 1
19787 kriscenter 1
19788 krisen 12
19789 krisens 1
19790 kriser 13
19791 krisförebyggande 1
19792 krisförordning 1
19793 krishantering 9
19794 krishanteringsplanerna 1
19795 krisläge 1
19796 krisläget 1
19797 krismedvetande 2
19798 krismöte 1
19799 krisområde 1
19800 krisområden 1
19801 krisperioden 1
19802 krisregionen 1
19803 krissituationen 1
19804 krissituationer 1
19805 krisstyrningsåtgärderna 1
19806 kristallklara 2
19807 kristdemokrater 20
19808 kristdemokraterna 5
19809 kristdemokraternas 1
19810 kristdemokratisk 1
19811 kristdemokratiska 1
19812 kristdemokratiske 1
19813 kristendom 1
19814 kristendomens 1
19815 kristna 1
19816 kritan 4
19817 kriterier 40
19818 kriterierna 8
19819 kriteriet 1
19820 kriterium 1
19821 kritik 28
19822 kritiken 10
19823 kritiker 2
19824 kritisera 18
19825 kritiserade 1
19826 kritiserades 1
19827 kritiserar 11
19828 kritiseras 3
19829 kritiserat 3
19830 kritiserats 1
19831 kritisk 20
19832 kritiska 17
19833 kritiskt 8
19834 kroater 1
19835 krocka 1
19836 krog 1
19837 krok 1
19838 krokar 2
19839 krokig 1
19840 krom 3
19841 krombrickor 1
19842 kromen 1
19843 kronan 1
19844 kronjuvelen 1
19845 kropp 9
19846 kroppar 3
19847 kroppen 4
19848 kroppens 1
19849 kropps 1
19850 kroppsbyggnad 1
19851 kroppslösa 1
19852 kroppsrytm 1
19853 kroppstemperatur 1
19854 krossa 1
19855 krossades 1
19856 krossar 1
19857 krukpalm 1
19858 krukskärva 1
19859 krumryggad 1
19860 krutdurk 1
19861 krutet 1
19862 krutröken 1
19863 kryddgården 1
19864 kryllar 1
19865 krympa 1
19866 krympande 1
19867 krypa 2
19868 kryphål 4
19869 kryphålen 1
19870 kryssa 1
19871 kryssningen 2
19872 kryssrutan 1
19873 kräftgång 1
19874 kränka 2
19875 kränkande 1
19876 kränker 5
19877 kränkning 9
19878 kränkningar 16
19879 kränkningarna 10
19880 kränks 5
19881 kränkt 1
19882 kränkta 1
19883 kränkts 1
19884 kräva 63
19885 krävande 7
19886 krävas 8
19887 krävde 6
19888 krävdes 7
19889 kräver 133
19890 krävs 147
19891 krävt 10
19892 krävts 2
19893 krångel 1
19894 krångla 1
19895 krånglar 1
19896 krånglig 1
19897 krångliga 1
19898 krökte 1
19899 krönas 1
19900 krönikör 2
19901 kröp 1
19902 kubanerna 1
19903 kubanernas 1
19904 kubansk 1
19905 kubanska 3
19906 kubikmeter 2
19907 kudde 1
19908 kudden 1
19909 kula 2
19910 kuliss 1
19911 kulisserna 4
19912 kullar 1
19913 kulle 1
19914 kullen 1
19915 kullerstensgatan 1
19916 kullerstensstenarna 1
19917 kullkasta 1
19918 kullkastar 1
19919 kullvräkt 1
19920 kulmen 1
19921 kulminerade 1
19922 kulor 1
19923 kulspetspenna 1
19924 kultiverad 1
19925 kultur 64
19926 kultur- 2
19927 kulturaktiviteter 1
19928 kulturanslag 1
19929 kulturarbetare 1
19930 kulturarv 7
19931 kulturarvet 2
19932 kulturell 19
19933 kulturella 26
19934 kulturella-historiska 1
19935 kulturellt 15
19936 kulturen 23
19937 kulturens 4
19938 kulturer 4
19939 kulturerna 1
19940 kulturform 1
19941 kulturförändring 1
19942 kulturhistoriskt 1
19943 kulturindustripolitik 1
19944 kulturområde 4
19945 kulturområdet 1
19946 kulturpolitik 5
19947 kulturpolitikens 1
19948 kulturpolitiska 1
19949 kulturprogram 2
19950 kulturprogrammet 1
19951 kulturresurserna 1
19952 kultursektorn 5
19953 kultursektors 1
19954 kulturservice 1
19955 kulturskillnader 1
19956 kulturutskottet 1
19957 kumulativa 3
19958 kumulativt 1
19959 kumuleringen 1
19960 kund 2
19961 kunde 237
19962 kunden 3
19963 kundens 1
19964 kunder 10
19965 kunderna 4
19966 kundernas 3
19967 kundkretsen 1
19968 kundorderformat 1
19969 kundorientering 1
19970 kundrelation 1
19971 kundvagnen 1
19972 kundvänliga 1
19973 kung 1
19974 kungariket 33
19975 kungarikets 12
19976 kungars 1
19977 kungen 1
19978 kungliga 1
19979 kungssportfiskare 1
19980 kunna 629
19981 kunnande 7
19982 kunnat 108
19983 kunnig 1
19984 kunnigt 1
19985 kunskap 26
19986 kunskapen 4
19987 kunskapens 2
19988 kunskaper 10
19989 kunskaperna 3
19990 kunskapsbaserad 3
19991 kunskapsbristen 1
19992 kunskapsdrivna 1
19993 kunskapsekonomi 2
19994 kunskapsekonomin 5
19995 kunskapsmässig 1
19996 kunskapsområdena 1
19997 kunskapssamhälle 4
19998 kunskapssamhället 7
19999 kunskapsspridning 1
20000 kunskapsträning 1
20001 kunskapsuppbyggnad 1
20002 kunskapsutveckling 1
20003 kunskapsöverföring 1
20004 kupolerna 1
20005 kurade 1
20006 kurder 1
20007 kurdiska 1
20008 kurs 5
20009 kursen 2
20010 kurser 1
20011 kurserna 1
20012 kursiv 1
20013 kursriktning 1
20014 kursändring 3
20015 kurva 2
20016 kusinen 1
20017 kusiner 1
20018 kuslig 2
20019 kusligt 1
20020 kust 7
20021 kust- 1
20022 kustbefolkningarnas 1
20023 kustbevakningen 1
20024 kustbevakningskårer 1
20025 kustbevakningsstyrka 1
20026 kusten 19
20027 kustens 2
20028 kuster 6
20029 kusterna 8
20030 kusternas 1
20031 kustfiskebåtar 1
20032 kustfisket 1
20033 kusthamnarna 1
20034 kustland 1
20035 kustlinje 2
20036 kustmyndigheter 2
20037 kustmyndigheternas 1
20038 kustneger 1
20039 kustnära 2
20040 kustområden 9
20041 kustområdena 3
20042 kustregioner 1
20043 kustregionerna 2
20044 kuststad 1
20045 kustvakter 1
20046 kustvatten 2
20047 kustvattnen 1
20048 kuvert 1
20049 kval 1
20050 kvalificera 2
20051 kvalificerad 20
20052 kvalificerade 8
20053 kvalificerat 3
20054 kvalifikationer 3
20055 kvalitativ 6
20056 kvalitativa 7
20057 kvalitativt 8
20058 kvalitet 55
20059 kvaliteten 34
20060 kvaliteter 2
20061 kvalitetsbevarande 1
20062 kvalitetsförbättringar 1
20063 kvalitetsförluster 1
20064 kvalitetsförsämring 1
20065 kvalitetsgaranti 1
20066 kvalitetskontroll 1
20067 kvalitetskrav 1
20068 kvalitetskraven 1
20069 kvalitetskriterier 1
20070 kvalitetsmärke 2
20071 kvalitetsmärkningens 1
20072 kvalitetsmätningen 1
20073 kvalitetsmålen 1
20074 kvalitetsnivå 1
20075 kvalitetsnormer 3
20076 kvalitetsprojekt 1
20077 kvalitetssprång 1
20078 kvalitetsvaror 1
20079 kvalitén 1
20080 kvalmigt 1
20081 kvantifierade 3
20082 kvantifieras 1
20083 kvantifierbara 4
20084 kvantitativ 3
20085 kvantitativa 9
20086 kvantitativt 3
20087 kvantitet 3
20088 kvantiteter 1
20089 kvantitetsgränser 1
20090 kvantitetshantering 1
20091 kvantitetshanteringen 1
20092 kvar 80
20093 kvarhängande 1
20094 kvarhålla 1
20095 kvarhållandena 1
20096 kvarhåller 1
20097 kvarhölls 1
20098 kvarleva 1
20099 kvarnsten 1
20100 kvarstad 1
20101 kvarstå 1
20102 kvarstår 10
20103 kvarstått 1
20104 kvartal 1
20105 kvartalet 1
20106 kvarter 8
20107 kvarteren 1
20108 kvarvarande 3
20109 kvasten 1
20110 kvastkäppen 1
20111 kvastskaft 1
20112 kvav 1
20113 kvavt 1
20114 kvestor 1
20115 kvestorer 3
20116 kvestorerna 9
20117 kvestorernas 1
20118 kvestorskollegiet 1
20119 kvickhet 1
20120 kvicksilver 6
20121 kvickt 1
20122 kvinna 31
20123 kvinnan 12
20124 kvinnans 4
20125 kvinnfolk 1
20126 kvinnlig 6
20127 kvinnliga 21
20128 kvinnlighet 1
20129 kvinnligt 2
20130 kvinnodagen 5
20131 kvinnofrågan 1
20132 kvinnogrupperna 1
20133 kvinnohandel 2
20134 kvinnokonferensen 1
20135 kvinnoprogrammet 2
20136 kvinnor 188
20137 kvinnorepresentationen 1
20138 kvinnorna 48
20139 kvinnornas 23
20140 kvinnors 45
20141 kvinnorörelsens 1
20142 kvinnoutskott 1
20143 kvinnoutskottet 1
20144 kvinnspersoner 1
20145 kvistar 1
20146 kvitt 2
20147 kvitterade 1
20148 kvot 10
20149 kvoten 3
20150 kvoter 17
20151 kvoterad 1
20152 kvotering 8
20153 kvoteringar 1
20154 kvoteringspolitik 1
20155 kvoteringspåföljder 1
20156 kvoterna 2
20157 kvotflyktingar 1
20158 kvotsystemet 1
20159 kväll 43
20160 kvällar 3
20161 kvällarna 2
20162 kvällen 13
20163 kvällens 4
20164 kvällningen 1
20165 kvällsflyget 1
20166 kvällsmat 1
20167 kvällsmöte 1
20168 kväva 4
20169 kväve 1
20170 kyckling 4
20171 kycklingar 2
20172 kycklingarna 1
20173 kycklingen 1
20174 kyla 3
20175 kylan 3
20176 kyliga 2
20177 kyligt 1
20178 kylskåpet 2
20179 kylstela 1
20180 kypare 1
20181 kyrka 1
20182 kyrkan 3
20183 kyrkans 2
20184 kyrkdörren 1
20185 kyrkogård 1
20186 kyrkorna 3
20187 kyrkpiano 1
20188 kyss 1
20189 kyssa 1
20190 kysste 1
20191 käbbel 1
20192 käbblade 1
20193 käckt 1
20194 käll- 1
20195 källa 15
20196 källan 5
20197 källare 1
20198 källaren 1
20199 källformat 1
20200 källor 8
20201 källorna 2
20202 kämpa 8
20203 kämpade 4
20204 kämpar 7
20205 kämpat 3
20206 känd 7
20207 kända 13
20208 kände 50
20209 kändes 15
20210 känga 1
20211 känn 2
20212 känna 41
20213 kännas 1
20214 kännbar 1
20215 kännbart 1
20216 kännedom 9
20217 kännedomen 1
20218 känner 170
20219 kännetecken 1
20220 känneteckna 2
20221 kännetecknade 1
20222 kännetecknades 2
20223 kännetecknande 1
20224 kännetecknar 1
20225 kännetecknas 7
20226 kännetecknat 1
20227 känns 3
20228 känsla 25
20229 känslan 13
20230 känslans 1
20231 känslig 23
20232 känsliga 17
20233 känsligare 2
20234 känsligaste 3
20235 känslighet 5
20236 känsligt 7
20237 känslokall 1
20238 känslokalla 1
20239 känsloladdad 1
20240 känslomässiga 2
20241 känslomässigt 1
20242 känslor 13
20243 känslotänkande 1
20244 känt 24
20245 känts 1
20246 käpp 1
20247 käpprakt 1
20248 kär 2
20249 kära 111
20250 käre 2
20251 kärl 2
20252 kärlek 6
20253 kärleken 4
20254 kärls 1
20255 kärna 6
20256 kärnaktivitet 1
20257 kärnan 8
20258 kärnenergisäkerhet 6
20259 kärnenergisäkerhetsfördragen 1
20260 kärnenergiäkerhet 1
20261 kärnfission 1
20262 kärnforskning 1
20263 kärnfrågan 2
20264 kärnfrågor 1
20265 kärnfusion 1
20266 kärnkatastrofer 1
20267 kärnkraft 5
20268 kärnkraften 1
20269 kärnkraftens 1
20270 kärnkraftsanläggningar 3
20271 kärnkraftsanläggningarna 1
20272 kärnkraftsolycka 1
20273 kärnkraftsolyckor 1
20274 kärnkraftsområdet 1
20275 kärnkraftsplanerna 1
20276 kärnkraftsprogram 1
20277 kärnkraftsreaktorer 1
20278 kärnkraftssäkerhet 1
20279 kärnkraftsverk 1
20280 kärnkraftverk 7
20281 kärnkraftverken 1
20282 kärnområden 1
20283 kärnprinciper 1
20284 kärnprinciperna 1
20285 kärnproblemen 1
20286 kärnpunkt 1
20287 kärnpunkten 2
20288 kärnpunkter 1
20289 kärnstrålningskontroller 1
20290 kärnsäkerhet 3
20291 kärnteknik 2
20292 kärnuppgifter 1
20293 kärnuppgifterna 1
20294 kärnvapen 6
20295 kärnvapenspridning 1
20296 kärnvapenteknik 1
20297 kärnvapenutveckling 1
20298 kärnverksamhet 1
20299 kärran 2
20300 kål 3
20301 kålhuven 1
20302 kånkande 1
20303 kår 1
20304 kåren 2
20305 kårer 1
20306 kåta 1
20307 kö 2
20308 köat 1
20309 köer 1
20310 kök 2
20311 köket 16
20312 köksbiträde 2
20313 köksbordet 3
20314 köksstol 1
20315 köksstolen 1
20316 köl 3
20317 kölar 1
20318 köld 3
20319 köldbeständigheten 1
20320 köldgränsen 1
20321 kölvattnet 1
20322 kön 12
20323 könen 15
20324 könens 1
20325 könet 1
20326 könsapartheid 1
20327 könsdiskriminering 1
20328 könsfrågor 1
20329 könsfördelning 2
20330 könsförändringar 1
20331 könsgrundade 1
20332 könsidentiteter 1
20333 könskvotering 5
20334 könsorgan 1
20335 könsrelaterad 1
20336 könsrelaterade 1
20337 könsspecifika 1
20338 köp 1
20339 köpa 5
20340 köpare 1
20341 köpas 1
20342 köpenskap 1
20343 köper 4
20344 köpet 4
20345 köpkraft 1
20346 köpkraften 1
20347 köpman 1
20348 köpmans 1
20349 köps 1
20350 köpslagningslogik 1
20351 köpslå 1
20352 köpt 4
20353 köpte 7
20354 kör 9
20355 köra 5
20356 köras 7
20357 körde 7
20358 kördes 1
20359 körförbud 1
20360 körning 1
20361 körningen 1
20362 körningsfel 1
20363 körs 3
20364 körsbärs- 1
20365 kört 4
20366 körtid 1
20367 körtidsfunktioner 1
20368 kött 2
20369 kött- 1
20370 köttkrig 1
20371 köttprodukter 1
20372 köttskiva 1
20373 l 1
20374 l'Etat 2
20375 l'Europe 1
20376 l'eau 1
20377 la 9
20378 laboratorier 1
20379 laboratorium 2
20380 laborerar 2
20381 labourkolleger 1
20382 labourledamöterna 1
20383 labourledamöternas 1
20384 labours 2
20385 labradoren 1
20386 labyrint 1
20387 lackerade 1
20388 lackstång 1
20389 lackstången 1
20390 laddat 2
20391 lade 53
20392 lades 18
20393 ladugårdsuggla 1
20394 lag 20
20395 laga 2
20396 lagade 2
20397 lagar 30
20398 lagarna 5
20399 lagbrott 1
20400 lagd 1
20401 lagen 19
20402 lagenligt 1
20403 lagens 2
20404 lager 6
20405 lagerhus 2
20406 lagerkrans 1
20407 laget 6
20408 lagförslag 6
20409 lagförslaget 2
20410 lagkränkning 1
20411 laglig 1
20412 lagliga 6
20413 laglighet 2
20414 lagligheten 1
20415 lagligt 8
20416 lagmängden 1
20417 lagom 1
20418 lagra 3
20419 lagrade 2
20420 lagrar 1
20421 lagras 1
20422 lagret 1
20423 lagring 1
20424 lagringskapacitet 1
20425 lags 1
20426 lagstadgad 1
20427 lagstadgade 2
20428 lagstifta 7
20429 lagstiftande 19
20430 lagstiftar 5
20431 lagstiftare 1
20432 lagstiftarna 2
20433 lagstiftat 2
20434 lagstiftning 125
20435 lagstiftningar 2
20436 lagstiftningen 59
20437 lagstiftningens 1
20438 lagstiftnings- 1
20439 lagstiftningsarbete 1
20440 lagstiftningsarbetet 6
20441 lagstiftningscykel 1
20442 lagstiftningsfrågor 1
20443 lagstiftningsförfarande 2
20444 lagstiftningsförfarandet 4
20445 lagstiftningsförslag 6
20446 lagstiftningsinitiativ 2
20447 lagstiftningsinstrument 1
20448 lagstiftningsmängd 1
20449 lagstiftningsområden 2
20450 lagstiftningsperioden 1
20451 lagstiftningsprocess 1
20452 lagstiftningsprocessen 5
20453 lagstiftningsprogram 9
20454 lagstiftningsprogrammet 8
20455 lagstiftningsprojektet 1
20456 lagstiftningsramen 1
20457 lagstiftningsreformen 1
20458 lagstiftningsresolutionen 10
20459 lagstiftningsresolutionerna 2
20460 lagstiftningsåtgärder 5
20461 lagt 105
20462 lagtext 2
20463 lagtexten 1
20464 lagtexter 1
20465 lagtexterna 1
20466 lagts 52
20467 lagändringar 1
20468 laissez 1
20469 lamaismen 1
20470 lambala-talande 1
20471 lamm 1
20472 lampa 1
20473 lampor 1
20474 lamporna 1
20475 lamslagen 1
20476 land 269
20477 landade 2
20478 landades 1
20479 landar 1
20480 landas 2
20481 landat 1
20482 landats 1
20483 landet 74
20484 landets 21
20485 landgränserna 2
20486 landminor 5
20487 landmärke 1
20488 landning 1
20489 landningen 2
20490 landningsbanan 1
20491 landområde 1
20492 landområden 1
20493 landpermission 2
20494 landremsan 1
20495 lands 15
20496 landsatte 3
20497 landsbruket 1
20498 landsbygd 3
20499 landsbygden 67
20500 landsbygdens 29
20501 landsbygdsbefolkningarna 1
20502 landsbygdsbefolkningen 1
20503 landsbygdskommuners 1
20504 landsbygdsområde 1
20505 landsbygdsområden 11
20506 landsbygdsområdena 3
20507 landsbygdsområdet 9
20508 landsbygdsområdets 1
20509 landsbygdspolitiken 1
20510 landsbygdsproblem 1
20511 landsbygdsregion 1
20512 landsbygdsregioner 2
20513 landsbygdsregionerna 2
20514 landsbygdsstrukturens 1
20515 landsbygdsturism 1
20516 landsbygdsutveckling 13
20517 landsbygdsutvecklingen 2
20518 landsbygdsutvecklingens 1
20519 landsflykten 1
20520 landsförvisning 2
20521 landskap 2
20522 landskapen 1
20523 landskapet 1
20524 landskapstrakter 1
20525 landsman 2
20526 landsmaninnor 2
20527 landsmän 6
20528 landsmäns 1
20529 landsspecifika 1
20530 landstiger 1
20531 landsväg 3
20532 landsändar 1
20533 landsätta 1
20534 landsättas 1
20535 landvinningar 4
20536 lansera 3
20537 lanserade 1
20538 lanserades 1
20539 lanserandet 1
20540 lanserar 1
20541 lanserat 1
20542 lansering 1
20543 lantbrukare 1
20544 lantbrukarna 1
20545 lantbruket 1
20546 lantbrukssamhälle 1
20547 lantdjur 1
20548 lantliga 1
20549 lappa 1
20550 lapptäcke 1
20551 lappverk 2
20552 larm 3
20553 larmrapporter 2
20554 larmsignal 2
20555 larver 1
20556 last 6
20557 lasta 2
20558 lastas 1
20559 lastat 1
20560 lastbalanserande 1
20561 lastbil 5
20562 lastbilar 6
20563 lastbilarna 2
20564 lastbilsförare 1
20565 lastbilskontroll 1
20566 lastbilsparken 1
20567 lastbilsstänkskärmar 1
20568 lastbilssäng 1
20569 lastbilsägare 1
20570 lastbilsägarna 1
20571 lasten 5
20572 lastens 2
20573 lasternas 1
20574 lastning 1
20575 lastområde 1
20576 lastrester 4
20577 lastrum 1
20578 lastångare 1
20579 latent 1
20580 latinamerikanska 1
20581 latituder 2
20582 latmansgöra 1
20583 lava 1
20584 law 2
20585 lax 7
20586 laxanemi 5
20587 laxanläggningar 1
20588 laxar 1
20589 laxen 2
20590 laxens 1
20591 laxindustrin 1
20592 laxodlare 1
20593 laxodlingar 1
20594 laxodlingsindustrin 1
20595 laxodlingssektorn 2
20596 laxrosa 1
20597 laxsektorn 1
20598 layout 6
20599 layouten 6
20600 le 6
20601 leasa 1
20602 led 4
20603 leda 122
20604 ledamot 99
20605 ledamoten 59
20606 ledamotens 6
20607 ledamotsstadga 1
20608 ledamotsstadgan 1
20609 ledamöter 159
20610 ledamöterna 58
20611 ledamöternas 9
20612 ledamöters 2
20613 ledande 15
20614 ledardjuren 1
20615 ledare 24
20616 ledaren 3
20617 ledarens 1
20618 ledares 1
20619 ledarförmåga 1
20620 ledarna 10
20621 ledarposition 1
20622 ledarskap 4
20623 ledarskapet 1
20624 ledas 2
20625 ledd 1
20626 ledda 2
20627 ledde 23
20628 leder 87
20629 ledet 3
20630 lediga 1
20631 ledmotiv 1
20632 ledning 16
20633 ledningar 1
20634 ledningen 14
20635 ledningscentralen 1
20636 ledningsförmågan 1
20637 ledningsmässiga 1
20638 ledningsnivåer 1
20639 ledningssätt 2
20640 ledningssättet 1
20641 ledningsutövning 1
20642 leds 2
20643 ledsaga 2
20644 ledsen 9
20645 ledstjärna 2
20646 ledstjärnan 1
20647 ledtrådar 1
20648 leende 18
20649 leendet 2
20650 legal 7
20651 legala 7
20652 legale 2
20653 legalisera 1
20654 legaliserade 1
20655 legalitet 5
20656 legaliteten 2
20657 legalitetsprincip 2
20658 legalt 9
20659 legat 5
20660 lege 1
20661 legender 1
20662 legionärerna 1
20663 legitim 3
20664 legitima 12
20665 legitimera 2
20666 legitimerar 2
20667 legitimeras 2
20668 legitimering 3
20669 legitimitet 10
20670 legitimiteten 3
20671 legitimt 1
20672 lejda 1
20673 lejer 1
20674 lejonporten 1
20675 leka 1
20676 lekarna 1
20677 lekbeståndens 1
20678 lekboll 1
20679 leker 3
20680 lekfullt 1
20681 lekområde 1
20682 lekplats 1
20683 leksaker 3
20684 lekt 1
20685 lekte 6
20686 lektion 1
20687 lektioner 3
20688 lektor 1
20689 lem 1
20690 lemlästande 1
20691 lemlästar 1
20692 lenande 1
20693 leninism 1
20694 leoparder 1
20695 ler 2
20696 lera 2
20697 leran 1
20698 lerhydda 1
20699 lerkärlen 1
20700 lerväggarna 1
20701 les 1
20702 leta 7
20703 letade 4
20704 letar 3
20705 letat 2
20706 lett 35
20707 leva 49
20708 levande 20
20709 levantinskt 1
20710 levat 1
20711 levde 8
20712 levebröd 5
20713 level 1
20714 lever 59
20715 leverans 1
20716 leveransen 1
20717 leverantör 1
20718 leverantörer 3
20719 leverantörskedjor 1
20720 leverar 1
20721 leverera 9
20722 levererar 2
20723 levereras 5
20724 levererat 3
20725 levnads- 1
20726 levnadsbetingelser 1
20727 levnadsglada 1
20728 levnadsnivå 1
20729 levnadsnivåer 1
20730 levnadsstandard 4
20731 levnadsstandarden 2
20732 levnadssätt 3
20733 levnadssättet 1
20734 levnadsvillkor 3
20735 levnadsvillkoren 1
20736 levt 3
20737 liaison 1
20738 libanesiska 2
20739 liberal 6
20740 liberala 56
20741 liberaldemokrater 1
20742 liberalen 1
20743 liberaler 3
20744 liberalerna 3
20745 liberalernas 1
20746 liberalisera 3
20747 liberalisering 4
20748 liberaliseringen 4
20749 liberalism 2
20750 liberalismen 2
20751 licens 1
20752 licenser 4
20753 licensfil 1
20754 licensiera 1
20755 licensinnehavarna 1
20756 licenspaketfil 1
20757 lida 6
20758 lidande 9
20759 lidanden 2
20760 lidandes 1
20761 lidandet 2
20762 lidelsefull 2
20763 lidelsefulla 4
20764 lider 21
20765 lidit 11
20766 lift 1
20767 liftare 1
20768 lifting 2
20769 liga 1
20770 ligga 34
20771 liggande 4
20772 ligger 184
20773 liggtidskostnaden 1
20774 lik 7
20775 lika 193
20776 likabehandling 1
20777 likaberättigad 1
20778 likadan 3
20779 likadana 3
20780 likadant 4
20781 likaledes 3
20782 likalydande 1
20783 likar 2
20784 likartad 1
20785 likartade 2
20786 likartat 1
20787 likaså 13
20788 likaväl 4
20789 likbleka 1
20790 likgiltig 2
20791 likgiltiga 4
20792 likgiltighet 2
20793 likgiltigheten 2
20794 likgiltigt 1
20795 likhet 34
20796 likheter 1
20797 likna 5
20798 liknade 7
20799 liknande 48
20800 liknar 14
20801 liknas 1
20802 liknat 1
20803 likriktade 4
20804 likriktande 1
20805 likriktas 1
20806 likriktning 2
20807 likriktningen 1
20808 liksidig 1
20809 liksom 158
20810 likstank 1
20811 likställa 3
20812 likställas 2
20813 likställda 2
20814 likställdes 1
20815 likställdhet 1
20816 likt 11
20817 likvida 2
20818 likväl 10
20819 likvärdig 4
20820 likvärdiga 8
20821 likvärdighet 1
20822 likvärdigt 1
20823 lila 1
20824 lilla 26
20825 lille 6
20826 lillfinger 2
20827 linan 1
20828 linbana 1
20829 linda 2
20830 lindra 4
20831 lindrande 1
20832 lindras 1
20833 lingua 1
20834 lingula 1
20835 lingvistiska 1
20836 linjal 1
20837 linjalen 1
20838 linjalens 1
20839 linje 35
20840 linjen 30
20841 linjer 5
20842 linjerna 4
20843 linjära 1
20844 linne 2
20845 linorna 1
20846 linsen 1
20847 lire 4
20848 lisa 1
20849 lista 13
20850 listan 13
20851 listigt 3
20852 listor 4
20853 listorna 2
20854 lita 6
20855 litade 2
20856 litar 10
20857 lite 36
20858 liten 73
20859 liter 1
20860 litet 147
20861 litteratur 7
20862 litteraturen 4
20863 litteraturförteckning 1
20864 litteraturförteckningen 1
20865 litterära 2
20866 liv 76
20867 livboj 1
20868 liverpoolskt 1
20869 livet 47
20870 livets 3
20871 livgardistuniform 1
20872 livlig 2
20873 livliga 5
20874 livligt 1
20875 livlina 2
20876 livnära 2
20877 livs 2
20878 livsbehov 2
20879 livsbesparingar 1
20880 livsbetingelserna 1
20881 livscykel 3
20882 livsdugliga 2
20883 livsförutsättningarna 1
20884 livshållning 1
20885 livskraft 2
20886 livskraften 1
20887 livskraftig 1
20888 livskraftiga 1
20889 livskvalitet 14
20890 livskvaliteten 9
20891 livskvalitén 2
20892 livslängden 1
20893 livslånga 1
20894 livslångt 9
20895 livsmedel 28
20896 livsmedels- 1
20897 livsmedelsbrist 2
20898 livsmedelsexport 1
20899 livsmedelsfrågor 1
20900 livsmedelsfrågorna 1
20901 livsmedelsföreskrifter 1
20902 livsmedelsföretagen 1
20903 livsmedelsförsörjningen 1
20904 livsmedelshanterares 1
20905 livsmedelshjälp 2
20906 livsmedelsindustrier 1
20907 livsmedelsindustrin 1
20908 livsmedelskedja 1
20909 livsmedelskedjan 2
20910 livsmedelskonsumtion 1
20911 livsmedelskontroll 2
20912 livsmedelskris 2
20913 livsmedelskriserna 1
20914 livsmedelskvalitet 3
20915 livsmedelslagstiftning 7
20916 livsmedelsmyndighet 8
20917 livsmedelsmyndigheten 4
20918 livsmedelsmyndighetens 1
20919 livsmedelsnyheterna 1
20920 livsmedelsområdet 1
20921 livsmedelsprodukter 1
20922 livsmedelsproduktion 1
20923 livsmedelsproduktionen 2
20924 livsmedelsproduktionskedjan 1
20925 livsmedelsprogram 1
20926 livsmedelssektorn 3
20927 livsmedelsstandarder 1
20928 livsmedelsstöd 1
20929 livsmedelssäkerhet 38
20930 livsmedelssäkerheten 7
20931 livsmedelssäkerhetens 1
20932 livsmedelssäkerhetsenheter 3
20933 livsmedelssäkerhetslagstiftningen 1
20934 livsmedelssäkerhetsmyndigheten 6
20935 livsmedelssäkerhetsmyndigheter 1
20936 livsmedelssäkerhetsområdet 1
20937 livsmedelssäkerhetssystem 1
20938 livsmedelstillverkningen 1
20939 livsmiljö 2
20940 livsmiljöer 6
20941 livsmiljöerna 1
20942 livsmiljön 1
20943 livsnödvändigt 1
20944 livspartner 1
20945 livsstil 1
20946 livstid 2
20947 livsuppehållande 1
20948 livsviktig 2
20949 livsviktigt 1
20950 livsvillkor 4
20951 livsyta 1
20952 livvakt 1
20953 ljud 11
20954 ljuda 1
20955 ljuder 1
20956 ljudet 4
20957 ljudlig 1
20958 ljudligt 1
20959 ljudlöst 1
20960 ljudupptagningar 6
20961 ljudupptagningar(11221/1999 1
20962 ljuga 2
20963 ljuger 1
20964 ljungeld 1
20965 ljus 20
20966 ljusa 8
20967 ljusan 1
20968 ljusare 2
20969 ljusblå 1
20970 ljusen 2
20971 ljuset 35
20972 ljushårig 1
20973 ljuskretsen 1
20974 ljuslagd 1
20975 ljuspunkter 1
20976 ljusrött 1
20977 ljussken 1
20978 ljusstråle 1
20979 ljustrafik 1
20980 ljusår 2
20981 ljuv 1
20982 ljuva 2
20983 ljuvlig 1
20984 ljuvliga 1
20985 ljuvligt 1
20986 lo 1
20987 lobby 1
20988 lobbyarbete 1
20989 lobbyarbetet 1
20990 lobbyföretag 1
20991 lobbygrupper 1
20992 lobbygrupperna 1
20993 lobbyintressen 1
20994 lobbymaskin 1
20995 lobbyverksamhet 3
20996 loca 1
20997 locka 4
20998 lockande 1
20999 lockar 1
21000 lockas 1
21001 lockats 1
21002 lockelse 2
21003 lockiga 1
21004 lockigt 2
21005 lodrät 1
21006 log 7
21007 loggade 1
21008 loggboken 1
21009 logik 9
21010 logiken 5
21011 logisk 1
21012 logiska 4
21013 logiskt 13
21014 logistik 2
21015 logistiken 1
21016 logistikorganisation 1
21017 logistikstöd 1
21018 loitering 1
21019 loj 1
21020 loja 1
21021 lojal 2
21022 lojalisterna 4
21023 lojalitet 1
21024 lojaliteten 1
21025 lojalt 3
21026 lojt 2
21027 lokal 27
21028 lokala 145
21029 lokalbefolkningen 3
21030 lokalen 1
21031 lokaler 4
21032 lokalerna 1
21033 lokaliseras 1
21034 lokalisering 2
21035 lokaliseringen 1
21036 lokaliseringsproblem 1
21037 lokalpatriotiska 1
21038 lokalpolis 1
21039 lokalsamhället 1
21040 lokalsamhällets 1
21041 lokalskatt 1
21042 lokalt 13
21043 lokaltidningen 1
21044 lokaltåg 1
21045 londonområdet 1
21046 look 1
21047 loopar 1
21048 lopp 9
21049 loppet 3
21050 loss 6
21051 lossa 1
21052 lossna 1
21053 lossnat 1
21054 lossning 1
21055 lots 1
21056 lotsade 1
21057 lotsat 1
21058 lotsens 1
21059 lotsning 1
21060 lott 2
21061 lottade 4
21062 lotusblomma 1
21063 lov 13
21064 lova 6
21065 lovade 19
21066 lovande 5
21067 lovar 7
21068 lovat 14
21069 lovats 1
21070 lovord 2
21071 lovorda 4
21072 lovordar 2
21073 lovordats 1
21074 lovprisar 1
21075 lovvärd 2
21076 lovvärda 3
21077 lovvärt 1
21078 lovyttringar 1
21079 lucka 4
21080 luckor 7
21081 luckorna 1
21082 luckra 1
21083 luddiga 3
21084 luddighet 1
21085 luddigt 2
21086 luft 7
21087 luftbro 1
21088 luftburet 1
21089 luftburna 1
21090 luften 21
21091 luftfarkost 1
21092 luftfart 1
21093 luftföroreningar 1
21094 luftkvalitet 1
21095 luftområde 1
21096 lufträder 1
21097 luftslottsbetänkande 1
21098 luftströmmarna 1
21099 lufttransport- 1
21100 lufttransporter 1
21101 lufttransporterna 1
21102 lugg 1
21103 luggar 1
21104 luggslitna 1
21105 lugn 11
21106 lugna 11
21107 lugnade 3
21108 lugnande 2
21109 lugnar 3
21110 lugnare 1
21111 lugnas 1
21112 lugne 1
21113 lugnt 6
21114 lukrativa 1
21115 lukt 1
21116 luktade 4
21117 luktar 1
21118 lukten 3
21119 lukter 1
21120 lumpsamlarverksamhet 1
21121 lunch 2
21122 lunchen 2
21123 luncher 1
21124 lunchtid 1
21125 lungor 1
21126 lur 1
21127 lura 1
21128 lurad 1
21129 lurande 1
21130 luras 3
21131 lurat 1
21132 luren 4
21133 lust 6
21134 lusten 1
21135 lustiga 3
21136 lustigare 1
21137 lustigt 1
21138 luta 2
21139 lutad 1
21140 lutade 12
21141 lutande 2
21142 lutar 1
21143 lutheranska 1
21144 lutning 1
21145 luxemburgare 1
21146 luxemburgska 1
21147 lycka 10
21148 lyckad 2
21149 lyckade 5
21150 lyckades 27
21151 lyckan 3
21152 lyckas 78
21153 lyckat 2
21154 lyckats 52
21155 lycklig 11
21156 lyckliga 4
21157 lyckligaste 1
21158 lyckligt 2
21159 lyckligtvis 6
21160 lyckojägare 1
21161 lyckosamt 2
21162 lycksalig 1
21163 lyckönska 7
21164 lyckönskas 1
21165 lyckönskningar 5
21166 lyckönskningsmeddelande 1
21167 lyda 4
21168 lydelse 4
21169 lyder 15
21170 lydigt 1
21171 lydnad 1
21172 lyft 3
21173 lyfta 20
21174 lyftade 1
21175 lyftas 1
21176 lyfte 9
21177 lyfter 3
21178 lyftkraftsteori 1
21179 lyhörd 1
21180 lyhördhet 2
21181 lykta 1
21182 lyktornas 1
21183 lynchad 1
21184 lynchningsscener 1
21185 lyrisk 1
21186 lyriska 1
21187 lysa 5
21188 lysande 11
21189 lyser 3
21190 lyssna 32
21191 lyssnade 17
21192 lyssnande 1
21193 lyssnar 14
21194 lyssnat 21
21195 lyssningsläge 1
21196 lyst 1
21197 lyste 4
21198 lyx 1
21199 lyxproblem 1
21200 läck 1
21201 läcka 2
21202 läckage 2
21203 läckan 1
21204 läckande 2
21205 läcker 4
21206 läckor 2
21207 läckt 4
21208 läckte 3
21209 läder 1
21210 läderaktigt 1
21211 läderpåse 1
21212 läge 29
21213 lägen 1
21214 lägena 1
21215 lägenhet 1
21216 lägenheten 8
21217 läger 2
21218 lägesbedömningar 1
21219 lägesrapport 2
21220 läget 24
21221 lägg 2
21222 lägga 216
21223 läggas 22
21224 lägger 76
21225 läggning 2
21226 läggs 46
21227 läglig 1
21228 lägliga 1
21229 lägligt 4
21230 lägre 27
21231 lägret 3
21232 lägst 2
21233 lägsta 7
21234 läkare 7
21235 läkaren 3
21236 läkarjobb 1
21237 läkarkontroller 2
21238 läkartjänst 1
21239 läkemedel 5
21240 läkemedelsindustrin 2
21241 läktarna 1
21242 läkte 1
21243 lämna 68
21244 lämnad 2
21245 lämnade 18
21246 lämnades 5
21247 lämnar 33
21248 lämnas 17
21249 lämnat 27
21250 lämnats 9
21251 lämningarna 1
21252 lämpa 1
21253 lämpad 1
21254 lämpade 3
21255 lämpar 2
21256 lämplig 27
21257 lämpliga 39
21258 lämpligare 4
21259 lämpligast 1
21260 lämpligaste 3
21261 lämpligen 1
21262 lämplighet 2
21263 lämpligheten 1
21264 lämplighetsprov 1
21265 lämpligt 67
21266 län 2
21267 länder 363
21268 länderna 135
21269 ländernas 18
21270 länders 14
21271 ländskynken 1
21272 längd 4
21273 längden 3
21274 länge 130
21275 längesedan 2
21276 längre 208
21277 längs 27
21278 längst 6
21279 längsta 1
21280 längtan 2
21281 längtar 3
21282 länk 10
21283 länka 3
21284 länkad 2
21285 länkade 1
21286 länken 1
21287 läppar 5
21288 läpparna 1
21289 läpparnas 1
21290 läppstift 1
21291 lär 7
21292 lära 35
21293 lärande 11
21294 lärandet 2
21295 lärare 4
21296 läraren 1
21297 lärarna 3
21298 läras 1
21299 lärd 1
21300 lärda 1
21301 lärde 7
21302 lärdom 13
21303 lärdomar 4
21304 lärjungar 1
21305 läroanstalter 1
21306 läroplanen 1
21307 lärorikt 1
21308 lärosatser 1
21309 lärs 1
21310 lärt 12
21311 lärts 1
21312 läs 3
21313 läsa 15
21314 läsare 2
21315 läsas 1
21316 läsbar 1
21317 läsbara 1
21318 läsbarare 1
21319 läser 24
21320 läsfrämjande 1
21321 läskunniga 1
21322 läskunnigheten 1
21323 läsmaterial 1
21324 läsning 1
21325 läsningen 1
21326 läst 16
21327 läste 16
21328 lät 17
21329 lätt 54
21330 lätta 8
21331 lättad 2
21332 lättade 1
21333 lättar 2
21334 lättare 39
21335 lättast 2
21336 lättaste 1
21337 lättat 1
21338 lättflytande 1
21339 lättförståelig 1
21340 lättförståeligt 1
21341 lätthet 1
21342 lättillgänglig 1
21343 lättillgängliga 1
21344 lättläst 1
21345 lättnad 4
21346 lättnader 3
21347 lättrogenhet 1
21348 lättsinnig 1
21349 lättsinnigt 1
21350 lättviktsfordon 1
21351 lättviktsmetoder 1
21352 lättvindigt 1
21353 lättvättat 1
21354 läxa 4
21355 läxan 3
21356 läxat 1
21357 läxor 4
21358 låda 2
21359 lådan 1
21360 lådfacks 1
21361 lådor 1
21362 lådorna 1
21363 låg 66
21364 låga 24
21365 låginkomsttagare 2
21366 låglönestrategierna 1
21367 lågorna 1
21368 lågt 9
21369 lån 4
21370 låna 1
21371 lånade 1
21372 lånat 1
21373 lånats 1
21374 lång 114
21375 lång- 1
21376 långa 56
21377 långdragen 2
21378 långdragna 1
21379 långfenad 1
21380 långfingret 1
21381 långfristig 1
21382 långfärdsbussar 1
21383 långrandig 2
21384 långrandigt 1
21385 långsam 1
21386 långsamhet 1
21387 långsamheten 1
21388 långsamma 6
21389 långsammare 3
21390 långsamt 25
21391 långsiktig 5
21392 långsiktiga 18
21393 långsiktighet 1
21394 långsiktigt 9
21395 långt 118
21396 långtgående 14
21397 långtids- 1
21398 långtidsarbetslösa 4
21399 långtidsarbetslöshet 5
21400 långtidsarbetslösheten 1
21401 långtifrån 3
21402 långtradare 2
21403 långvariga 8
21404 långvarigt 4
21405 lår 1
21406 låsa 4
21407 låser 2
21408 låset 1
21409 låsningarna 1
21410 låsningen 1
21411 låst 2
21412 låsta 1
21413 låsts 1
21414 låt 47
21415 låta 106
21416 låter 33
21417 låtit 6
21418 låtsad 1
21419 låtsades 1
21420 låtsas 10
21421 löddrade 1
21422 löfte 14
21423 löften 21
21424 löftena 1
21425 löftesrika 1
21426 löftesrikt 1
21427 löftet 4
21428 lögn 1
21429 lögnen 1
21430 lögner 2
21431 löjeväckande 4
21432 löjlig 1
21433 löjliga 1
21434 löjligt 1
21435 lökar 1
21436 lökformade 2
21437 lökmodell 1
21438 lömsk 1
21439 lömskt 1
21440 lön 8
21441 löna 2
21442 lönar 1
21443 löne- 3
21444 lönearbetsrättigheter 1
21445 lönebesked 2
21446 löneeffektivitet 1
21447 löneförhållandena 1
21448 lönehöjningarna 1
21449 lönemässigt 1
21450 lönen 2
21451 lönepaketet 1
21452 lönepolitik 3
21453 löner 8
21454 lönerna 2
21455 lönetak 1
21456 löneökningar 1
21457 löneökningspolitik 1
21458 lönsam 3
21459 lönsamhet 2
21460 lönsamhets- 1
21461 lönsamhetstänkande 1
21462 lönsamma 6
21463 lönsamt 2
21464 lönt 2
21465 löntagare 2
21466 löntagarna 6
21467 löpa 4
21468 löpande 11
21469 löpeld 1
21470 löper 13
21471 löpt 6
21472 löpte 5
21473 lördag 3
21474 lördagskvällar 1
21475 lös 7
21476 lösa 103
21477 lösare 1
21478 lösas 16
21479 lösenord 1
21480 lösenordet 3
21481 löser 10
21482 löses 2
21483 lösesumma 1
21484 lösgör 1
21485 lösning 109
21486 lösningar 52
21487 lösningarna 1
21488 lösningen 23
21489 lösningsförslag 1
21490 lösnäsa 1
21491 lösryckt 1
21492 löst 10
21493 lösta 5
21494 löste 2
21495 löstes 3
21496 lösts 9
21497 löv 1
21498 löven 1
21499 lövskogarna 1
21500 m 1
21501 m.fl. 3
21502 m.m. 5
21503 m3 2
21504 mader 1
21505 maffia 1
21506 maffian 1
21507 maffians 1
21508 maffior 1
21509 magasin 3
21510 magasinerade 2
21511 mage 3
21512 magen 5
21513 mager 5
21514 magi 4
21515 magisk 2
21516 magiska 3
21517 magiskt 1
21518 magknipande 2
21519 magnet 1
21520 magnifik 1
21521 magnifika 1
21522 magnitud 1
21523 magra 1
21524 magrare 1
21525 magstarkt 1
21526 mainstraming 1
21527 mainstreaming 18
21528 mainstreaming-program 1
21529 maj 23
21530 majestätiskt 1
21531 majoritet 54
21532 majoriteten 19
21533 majoriteter 1
21534 majoriteterna 1
21535 majoritetsbeslut 4
21536 majoritetsbeslutet 1
21537 majoritetsgrupp 1
21538 majoritetsomröstningar 1
21539 majoritetsröstning 1
21540 majoritetsuppfattning 1
21541 majoritetsuppfattningen 1
21542 majs 1
21543 makabert 1
21544 makade 1
21545 makarna 2
21546 make 2
21547 makedonierna 3
21548 makedonisk 1
21549 makedoniska 7
21550 makedoniskt 1
21551 maken 1
21552 makroekonomin 1
21553 makroekonomisk 5
21554 makroekonomiska 17
21555 makroekonomiskt 3
21556 makrofinansiellt 1
21557 makropolitik 1
21558 makt 40
21559 maktambitioner 1
21560 maktbalans 1
21561 maktbalansen 1
21562 maktbefogenhet 3
21563 maktbefogenheter 2
21564 maktberusning 1
21565 maktcentrumen 1
21566 maktdelningen 1
21567 maktdikterade 1
21568 makten 23
21569 maktens 2
21570 makter 2
21571 makterna 1
21572 maktfaktor 2
21573 maktförlusten 1
21574 makthavare 2
21575 makthavarna 2
21576 maktkoncentration 2
21577 maktkoncentrationen 1
21578 maktkoncentrationer 1
21579 maktlös 4
21580 maktlösa 1
21581 maktlöshet 3
21582 maktlöst 1
21583 maktmedel 3
21584 maktmedlen 1
21585 maktmissbruk 3
21586 maktpolitiska 1
21587 maktpositionen 1
21588 maktpositioner 2
21589 maktstrukturer 1
21590 maktövertagande 1
21591 mal 1
21592 malaria 1
21593 malariamyggan 1
21594 maldes 1
21595 mall 3
21596 malplacerade 1
21597 malt 1
21598 maltesarna 1
21599 malteserna 1
21600 maltesisk 3
21601 maltesiska 2
21602 maltwhisky 1
21603 maltwhiskyproducerande 1
21604 malört 1
21605 mamma 8
21606 mammas 1
21607 man 1905
21608 mana 2
21609 manad 1
21610 manade 1
21611 management 1
21612 managementnivå 1
21613 manar 4
21614 manas 1
21615 manat 1
21616 mandat 20
21617 mandaten 1
21618 mandatet 4
21619 mandatperiod 15
21620 mandatperioden 10
21621 mandatperiodens 2
21622 mandel 1
21623 maner 1
21624 mangoträden 1
21625 mangoträdens 1
21626 mangroveträden 1
21627 manifestationen 1
21628 manifestationer 1
21629 manifestationerna 1
21630 manifesterar 1
21631 maning 2
21632 manipulation 2
21633 manipulerad 1
21634 manlig 2
21635 manliga 11
21636 manligt 1
21637 manna 1
21638 mannen 26
21639 mannens 2
21640 mans 1
21641 manschetter 1
21642 manschettknappar 1
21643 manteln 1
21644 mantra 1
21645 mantran 1
21646 mantrat 1
21647 manuella 1
21648 manuellt 1
21649 manuskript 1
21650 manuskriptet 1
21651 manuskriptsamling 1
21652 manér 1
21653 manöver 2
21654 manövern 1
21655 manövrer 1
21656 manövrerade 1
21657 mapp 1
21658 mapparna 2
21659 mappen 2
21660 maratonlångt 1
21661 mardröm 1
21662 mardrömmar 3
21663 mardrömslik 1
21664 marginal 3
21665 marginalen 4
21666 marginaler 3
21667 marginalerna 1
21668 marginalisera 3
21669 marginaliserade 5
21670 marginaliserats 1
21671 marginalisering 2
21672 marginellt 2
21673 marin 2
21674 marina 18
21675 marionett 1
21676 maris 2
21677 maritima 2
21678 maritimt 2
21679 mark 13
21680 markant 4
21681 markanta 1
21682 markanvändning 1
21683 marken 13
21684 markens 1
21685 markera 2
21686 markerad 3
21687 markerade 2
21688 markerades 1
21689 markerar 10
21690 markeras 2
21691 markerat 2
21692 markering 3
21693 market 1
21694 marknad 50
21695 marknaden 192
21696 marknadens 26
21697 marknader 21
21698 marknaderna 18
21699 marknadernas 7
21700 marknadsaktören 1
21701 marknadsaktörerna 1
21702 marknadsaktörernas 1
21703 marknadsandel 2
21704 marknadsandelar 8
21705 marknadsdominans 1
21706 marknadsekonomi 13
21707 marknadsekonomin 8
21708 marknadsekonomins 2
21709 marknadsekonomiska 3
21710 marknadsföring 2
21711 marknadsföringskoncept 1
21712 marknadsinstrumentet 1
21713 marknadskrafter 1
21714 marknadskrafterna 1
21715 marknadslagarna 1
21716 marknadsliberalism 1
21717 marknadsmöjlighet 1
21718 marknadsorganisation 1
21719 marknadsorganisationen 1
21720 marknadspriser 2
21721 marknadsproblem 2
21722 marknadsprodukt 1
21723 marknadssituation 1
21724 marknadstillträde 4
21725 marktrupper 1
21726 marmorbyggnad 1
21727 marmortrappan 1
21728 marockanska 4
21729 marokäng 1
21730 mars 56
21731 marschera 1
21732 marscherande 1
21733 marscherar 1
21734 marshmallow 1
21735 marshmallow-klunsar 1
21736 marshmallowen 1
21737 marshmallows 1
21738 marskalken 1
21739 marskgräs 1
21740 marskgräset 2
21741 martinis 1
21742 mask 2
21743 masker 1
21744 maskerad 1
21745 maskin 3
21746 maskinellt 1
21747 maskinen 2
21748 maskiner 1
21749 maskineri 2
21750 maskineriet 2
21751 maskinist 1
21752 maskinistexamen 1
21753 maskinrummen 1
21754 maskinrummet 1
21755 maskinskada 1
21756 maskopi 1
21757 maskstungna 1
21758 masochister 1
21759 masochistisk 1
21760 masochistiska 1
21761 massa 11
21762 massaker 1
21763 massakerplatserna 1
21764 massakrera 1
21765 massakrerade 1
21766 massakrerna 1
21767 massan 1
21768 massans 1
21769 massarbetslöshet 1
21770 massarbetslösheten 2
21771 massavgång 1
21772 massiv 3
21773 massiva 7
21774 massivt 2
21775 massmedia 4
21776 massmedias 2
21777 massorna 1
21778 massrörelse 1
21779 masten 1
21780 masterna 1
21781 mastodont 1
21782 mat 13
21783 mata 1
21784 matade 1
21785 matat 1
21786 matbricka 1
21787 match 3
21788 matcha 2
21789 matchande 1
21790 matchar 2
21791 matdags 1
21792 matematiker 1
21793 matematisk 1
21794 matematiska 1
21795 maten 3
21796 material 28
21797 materialanskaffning 1
21798 materialen 1
21799 materialet 3
21800 materiell 1
21801 materiella 2
21802 materiellt 2
21803 matlagning 1
21804 matnyttiga 1
21805 matpaket 2
21806 matpensioner 1
21807 matrester 1
21808 matroserna 1
21809 matsal 1
21810 matsalen 3
21811 matsalsfönstret 1
21812 matsedeln 1
21813 matsedlarna 1
21814 matstrupe 1
21815 matt 1
21816 matta 1
21817 mattan 3
21818 mattorna 1
21819 maxbeloppen 1
21820 maximal 7
21821 maximala 3
21822 maximalt 7
21823 maximera 4
21824 maximerar 1
21825 maximistraffet 1
21826 maxstraffet 1
21827 maxvikter 1
21828 med 5242
21829 medaljbehängda 1
21830 medan 115
21831 medansvar 3
21832 medarbetare 7
21833 medbeslutande 14
21834 medbeslutandeförfarande 3
21835 medbeslutandeförfarandet 11
21836 medbeslutanderätt 3
21837 medbeslutandet 3
21838 medborgardebatt 1
21839 medborgardebatter 1
21840 medborgardemonstration 1
21841 medborgare 142
21842 medborgaren 21
21843 medborgaren-konsumenten 1
21844 medborgarens 1
21845 medborgares 18
21846 medborgarna 170
21847 medborgarnas 59
21848 medborgarrätt 1
21849 medborgarrörelser 1
21850 medborgarsamhället 2
21851 medborgarskap 6
21852 medborgarskapet 4
21853 medborgarskapsbegrepp 1
21854 medborgarskapsregleringen 1
21855 medborgarstadga 1
21856 medborgartanken 1
21857 medborgarvärde 1
21858 medborgerlig 1
21859 medborgerliga 21
21860 medborgerligt 2
21861 medbroders 1
21862 medbrottslighet 1
21863 medbrottslingar 1
21864 meddela 25
21865 meddelade 7
21866 meddelades 1
21867 meddelande 89
21868 meddelanden 12
21869 meddelandeskyldigheten 1
21870 meddelandet 34
21871 meddelandetexten 1
21872 meddelar 7
21873 meddelat 5
21874 medel 165
21875 medel- 1
21876 medelklass 3
21877 medellängd 1
21878 medellång 13
21879 medelmåttan 1
21880 medelmåttiga 1
21881 medelpunkt 2
21882 medelst 1
21883 medelstor 3
21884 medelstora 72
21885 medelstort 1
21886 medeltida 3
21887 medeltiden 1
21888 medelvärden 1
21889 medelålder 1
21890 medelåldern 1
21891 medelålders 3
21892 medfarna 1
21893 medfinansierade 1
21894 medfinansieras 1
21895 medfinansiering 1
21896 medfinansieringen 1
21897 medföljde 1
21898 medför 44
21899 medföra 17
21900 medförde 3
21901 medföredragande 2
21902 medfört 5
21903 medgav 2
21904 medge 7
21905 medger 24
21906 medges 9
21907 medgett 1
21908 medgivande 2
21909 medgivits 2
21910 medgörliga 1
21911 medgörlighet 1
21912 medhjälpare 1
21913 media 11
21914 mediaföretagen 1
21915 medial 1
21916 mediatäckningen 1
21917 medicin 2
21918 mediciner 1
21919 medicinsk 3
21920 medicinska 1
21921 medie- 1
21922 medier 7
21923 medierna 4
21924 mediernas 3
21925 medinflytande 2
21926 meditera 1
21927 medkänsla 9
21928 medla 2
21929 medlare 1
21930 medlaren 1
21931 medlem 25
21932 medlemmar 42
21933 medlemmarna 2
21934 medlemmars 1
21935 medlemsavgifter 1
21936 medlemskandidaterna 1
21937 medlemskap 23
21938 medlemskapet 1
21939 medlemskapsförhandlingarna 4
21940 medlemskapsprocessen 2
21941 medlemskapsrättigheter 1
21942 medlemskapsstöden 1
21943 medlemskapsåtgärder 1
21944 medlemsland 12
21945 medlemslandet 3
21946 medlemslands 1
21947 medlemsländer 21
21948 medlemsländerna 38
21949 medlemsländernas 12
21950 medlemsländers 2
21951 medlemsregeringarnas 1
21952 medlemsstarter 1
21953 medlemsstat 88
21954 medlemsstaten 15
21955 medlemsstatens 3
21956 medlemsstater 196
21957 medlemsstaterna 330
21958 medlemsstaterna- 1
21959 medlemsstaternas 90
21960 medlemsstaters 9
21961 medlemsstats 13
21962 medlemsstatsnivå 7
21963 medlemsstatsrapport 1
21964 medlen 20
21965 medlet 2
21966 medlidande 2
21967 medling 1
21968 medlingsförfarande 3
21969 medlingsförsök 1
21970 medlingsförsöken 1
21971 medlingsprocess 1
21972 medmänniskor 1
21973 medmänniskors 1
21974 medmänskliga 1
21975 medmänsklighet 2
21976 medskyldiga 2
21977 medspelarna 1
21978 medsvuren 1
21979 medverka 17
21980 medverkade 1
21981 medverkan 12
21982 medverkar 9
21983 medverkat 4
21984 medvetande 9
21985 medvetandehöjande 1
21986 medvetandenivå 1
21987 medvetandet 1
21988 medveten 47
21989 medvetenhet 7
21990 medvetenheten 1
21991 medvetet 13
21992 medvetna 60
21993 medvetslöshet 1
21994 megaprojekt 1
21995 mej 1
21996 mejeriindustrin 1
21997 meka 1
21998 mekanik 1
21999 mekanisk 2
22000 mekaniska 3
22001 mekaniskt 3
22002 mekanism 5
22003 mekanismen 1
22004 mekanismer 18
22005 mekanismerna 7
22006 mekanistiska 1
22007 mellan 738
22008 mellanfolklig 1
22009 mellanlagras 1
22010 mellanlagringar 1
22011 mellanled 2
22012 mellanliggande 5
22013 mellannivå 1
22014 mellanrum 1
22015 mellanskillnaden 1
22016 mellanstadiet 1
22017 mellanstatlig 5
22018 mellanstatliga 2
22019 mellanstatligt 6
22020 mellanstora 2
22021 mellanting 1
22022 mellanvägg 1
22023 mellanöstern 1
22024 membre 2
22025 memoarer 1
22026 men 1351
22027 mena 1
22028 menade 13
22029 menar 70
22030 menas 3
22031 mening 93
22032 meningar 3
22033 meningarna 1
22034 meningen 16
22035 meningsfull 4
22036 meningsfulla 3
22037 meningsfullt 14
22038 meningslös 4
22039 meningslösa 2
22040 meningslöst 7
22041 meningsskiljaktigheter 8
22042 meningsskiljaktigheterna 1
22043 menligt 1
22044 mentala 1
22045 mentalitet 1
22046 mentaliteten 5
22047 mentalsjuk 1
22048 meny 1
22049 menyn 3
22050 mer 619
22051 mera 60
22052 merger 1
22053 meriter 4
22054 meritokrati 1
22055 merkostnaden 1
22056 merparten 1
22057 mervärde 10
22058 mervärdesskattesats 1
22059 mervärdesstruktur 1
22060 mervärdet 1
22061 mesanmasten 1
22062 mest 149
22063 mesta 11
22064 mestadels 2
22065 metaforen 1
22066 metafysiskt 1
22067 metall 1
22068 metaller 3
22069 metallindustrin 1
22070 metalliska 1
22071 meter 4
22072 metersystemet 1
22073 metervis 1
22074 metod 29
22075 metoden 9
22076 metoder 36
22077 metoderna 5
22078 metodik 1
22079 metodiken 3
22080 metodikens 1
22081 metodikändringar 1
22082 metodiskt 4
22083 metodutveckling 1
22084 middag 4
22085 middagen 6
22086 middagsbjudningen 1
22087 middagsbord 1
22088 middagsbordet 1
22089 middagsgäster 1
22090 middagsgästerna 1
22091 middagshetta 1
22092 midja 1
22093 midjan 2
22094 midnatt 2
22095 mig 798
22096 migration 2
22097 migrationen 2
22098 migrationsrörelser 1
22099 migrationsströmmar 2
22100 migrationsströmmen 1
22101 mikrober 1
22102 mikroföretag 2
22103 mikrokrediter 2
22104 mikroprojekt 1
22105 mikrostater 1
22106 mikrostaterna 1
22107 mild 2
22108 mildare 1
22109 mildaste 1
22110 mildra 8
22111 mildrande 1
22112 mildras 1
22113 milen 1
22114 milis 2
22115 militariserade 1
22116 militarisering 2
22117 militarismen 1
22118 militär 20
22119 militära 52
22120 militäraktion 1
22121 militäraktioner 1
22122 militärer 2
22123 militärerna 1
22124 militärindustri 1
22125 militärinsats 1
22126 militärinsatserna 1
22127 militärkupp 1
22128 militärläger 1
22129 militärpolitiken 1
22130 militärsamarbete 1
22131 militärstyrkorna 1
22132 militärstyrkornas 1
22133 militärt 4
22134 militäruniformer 1
22135 miljard 1
22136 miljarder 40
22137 miljon 10
22138 miljoner 176
22139 miljonerna 3
22140 miljontals 3
22141 miljö 98
22142 miljö- 8
22143 miljöanpassad 2
22144 miljöansvar 3
22145 miljöansvaret 2
22146 miljöansvariga 1
22147 miljöarbete 1
22148 miljöarbetet 3
22149 miljöaspekten 4
22150 miljöaspekter 1
22151 miljöaspekterna 5
22152 miljöavtal 1
22153 miljöbelastningen 1
22154 miljöberoendet 1
22155 miljöbeskattning 1
22156 miljöbeskattningen 1
22157 miljöbestämmelser 1
22158 miljöbestämmelserna 1
22159 miljöbovar 1
22160 miljöbovarna 1
22161 miljöbrott 1
22162 miljöbrottsmyndighet 1
22163 miljöcowboys 1
22164 miljödepartementet 1
22165 miljödimensionen 2
22166 miljödirektiv 3
22167 miljödirektiven 1
22168 miljödirektivet 1
22169 miljödirektoratet 1
22170 miljödogmatism 1
22171 miljöeffekter 1
22172 miljöer 5
22173 miljöexperter 1
22174 miljöfaktor 1
22175 miljöfarliga 1
22176 miljöfråga 1
22177 miljöfrågan 1
22178 miljöfrågor 11
22179 miljöfrågorna 3
22180 miljöförbättrande 1
22181 miljöförbättring 1
22182 miljöfördelar 1
22183 miljöförhållandena 1
22184 miljöförordningen 1
22185 miljöförstörande 1
22186 miljöförstörelse 2
22187 miljöförstöring 5
22188 miljöförstöringen 1
22189 miljöförsämring 1
22190 miljögrupper 1
22191 miljöhänsyn 10
22192 miljöhänsynen 1
22193 miljöinformation 1
22194 miljöinsatserna 1
22195 miljökastastrofen 1
22196 miljökatastrof 12
22197 miljökatastrofala 1
22198 miljökatastrofen 3
22199 miljökatastrofens 1
22200 miljökatastroferna 1
22201 miljökommissionär 1
22202 miljökommissionären 1
22203 miljökonferensen 1
22204 miljökonsekvensbedömning 2
22205 miljökonsekvensbeskrivning 1
22206 miljökonsekvenser 5
22207 miljökonsekvenserna 3
22208 miljökostnaderna 2
22209 miljökrav 6
22210 miljökraven 4
22211 miljökriterierna 1
22212 miljökunskap 1
22213 miljökvaliteten 1
22214 miljölagstiftning 3
22215 miljölagstiftningen 2
22216 miljölagstiftningens 1
22217 miljömedvetandet 2
22218 miljömetoder 1
22219 miljöminister 3
22220 miljöministern 1
22221 miljöministrarna 1
22222 miljömyndigheterna 1
22223 miljömässig 2
22224 miljömässiga 18
22225 miljömässigt 5
22226 miljömål 5
22227 miljömålen 1
22228 miljömålsättningarna 1
22229 miljön 123
22230 miljönormer 2
22231 miljönormerna 2
22232 miljöns 3
22233 miljönätverk 1
22234 miljöområde 1
22235 miljöområden 2
22236 miljöområdet 13
22237 miljöorgan 1
22238 miljöorganisation 1
22239 miljöovänligt 1
22240 miljöpartist 1
22241 miljöpelaren 1
22242 miljöperspektiv 1
22243 miljöpolicyavtal 1
22244 miljöpolitik 7
22245 miljöpolitiken 7
22246 miljöpolitikens 1
22247 miljöpolitisk 1
22248 miljöpolitiska 2
22249 miljöpolitiskt 3
22250 miljöproblem 5
22251 miljöproblemen 3
22252 miljöprogram 1
22253 miljöprogrammen 1
22254 miljöprogrammering 1
22255 miljöprojekt 1
22256 miljöpåverkan 4
22257 miljöregelverket 1
22258 miljörelaterade 1
22259 miljöresultat 1
22260 miljörisker 1
22261 miljörådet 1
22262 miljörörelsen 3
22263 miljörörelsens 1
22264 miljörörelserna 1
22265 miljösektorerna 1
22266 miljösidan 1
22267 miljösituationen 1
22268 miljöskadliga 2
22269 miljöskador 2
22270 miljöskydd 16
22271 miljöskyddet 5
22272 miljöskyddets 1
22273 miljöskyddsbehoven 1
22274 miljöskyddsnivå 2
22275 miljöskyddsområdet 1
22276 miljöskyddspolitik 1
22277 miljöskyddsstöd 1
22278 miljöskäl 3
22279 miljöstudier 1
22280 miljöstöd 1
22281 miljösyften 1
22282 miljösynpunkt 8
22283 miljötragedi 1
22284 miljötvånget 1
22285 miljöuppgifter 2
22286 miljöutskottet 7
22287 miljöutskottets 1
22288 miljövariabler 1
22289 miljövänlig 2
22290 miljövänliga 7
22291 miljövänligaste 1
22292 miljövänligt 4
22293 miljövärdena 2
22294 miljöövervakningsenhet 1
22295 milkshakes 1
22296 millenniefebern 1
22297 millenniefusioner 1
22298 millennieskifte 1
22299 millennieskiftet 2
22300 millenniet 4
22301 millennietal 1
22302 millenniets 1
22303 millennium 2
22304 millimeteranpassade 1
22305 milstolpar 1
22306 milstolpe 3
22307 min 518
22308 min. 2
22309 mina 214
22310 minamatasjukdomen 1
22311 mindervärdiga 1
22312 minderårig 1
22313 minderåriga 3
22314 mindes 3
22315 mindre 184
22316 minen 1
22317 mineraler 1
22318 miniatyr 2
22319 minimal 1
22320 minimala 1
22321 minimalistiska 1
22322 minimalistiskt 1
22323 minimera 6
22324 minimeras 1
22325 minimibelopp 1
22326 minimibestämmelser 2
22327 minimifinansiering 1
22328 minimigemenskapsprogram 1
22329 minimiinkomst 1
22330 minimiinnehållet 1
22331 minimiinsatser 1
22332 minimikalender 1
22333 minimikapital 1
22334 minimikontroll 1
22335 minimikrav 4
22336 minimikraven 1
22337 minimikvoter 1
22338 minimilängden 1
22339 minimilön 1
22340 minimilönen 1
22341 minimilöner 2
22342 miniminivå 2
22343 miniminivån 1
22344 miniminormer 5
22345 minimipensionerna 1
22346 minimiprogram 1
22347 minimiprogrammet 2
22348 minimireform 2
22349 minimireformer 1
22350 minimiregler 5
22351 minimireglerna 2
22352 minimirättigheterna 1
22353 minimis-notis 1
22354 minimiskatter 1
22355 minimistandarden 1
22356 minimistandarder 2
22357 minimitaket 1
22358 minimitarifferna 1
22359 minimiuppehälle 1
22360 minimivikt 1
22361 minimiåtgärder 1
22362 minimorum 1
22363 minimum 12
22364 minireform 1
22365 minister 17
22366 ministerier 1
22367 ministermöte 1
22368 ministermötet 3
22369 ministern 16
22370 ministernivå 1
22371 ministerns 1
22372 ministerpost 1
22373 ministerposter 2
22374 ministerpresidenten 3
22375 ministerråd 5
22376 ministerrådet 22
22377 ministerrådets 1
22378 ministerrådsmöte 1
22379 ministrar 16
22380 ministrarna 8
22381 ministrars 1
22382 mink 1
22383 minkpäls 1
22384 minnas 6
22385 minne 11
22386 minnen 2
22387 minnena 2
22388 minnens 1
22389 minnesbild 1
22390 minnesmärke 1
22391 minnestal 1
22392 minnesvärda 1
22393 minnet 9
22394 minns 23
22395 minore 1
22396 minoritet 16
22397 minoriteten 7
22398 minoritetens 1
22399 minoriteter 25
22400 minoriteterna 6
22401 minoriteternas 2
22402 minoriteters 2
22403 minoritetsbefolkningar 1
22404 minoritetsfientliga 1
22405 minoritetsgrupper 5
22406 minoritetspolitik 1
22407 minoritetspolitiken 1
22408 minoritetsregering 3
22409 minorna 1
22410 minpolitiken 1
22411 minröjning 1
22412 minsann 2
22413 minska 87
22414 minskad 13
22415 minskade 11
22416 minskades 2
22417 minskande 4
22418 minskar 26
22419 minskas 9
22420 minskat 17
22421 minskats 2
22422 minskning 38
22423 minskningar 3
22424 minskningen 8
22425 minst 98
22426 minsta 31
22427 minste 1
22428 minttabletter 1
22429 minus 3
22430 minusgrader 2
22431 minut 13
22432 minuten 2
22433 minuter 24
22434 minuters 1
22435 minåtgärdsprogrammens 1
22436 mirakel 2
22437 mirakellösning 1
22438 mirakelmedel 1
22439 mirakulöst 1
22440 missa 3
22441 missade 2
22442 missat 4
22443 missbelåtenhet 1
22444 missbruk 14
22445 missbruka 1
22446 missbrukade 1
22447 missbrukades 1
22448 missbrukar 1
22449 missbrukas 1
22450 missbrukat 1
22451 missbruket 2
22452 missbruksprincipen 1
22453 missfall 1
22454 missfallen 2
22455 missfoster 1
22456 missförhållande 2
22457 missförhållandena 1
22458 missförhållandet 1
22459 missförstod 2
22460 missförstå 1
22461 missförstånd 7
22462 missförstår 1
22463 missförstås 1
22464 missgynna 2
22465 missgynnade 14
22466 missgynnas 1
22467 misshandel 3
22468 misshandlade 1
22469 misshandlar 1
22470 misshushållning 2
22471 mission 2
22472 missions 1
22473 missionsskolan 1
22474 missionären 1
22475 misskreditera 1
22476 misskrediterar 1
22477 misskötsel 7
22478 misskött 1
22479 misslyckad 1
22480 misslyckade 5
22481 misslyckades 5
22482 misslyckande 14
22483 misslyckanden 5
22484 misslyckandet 2
22485 misslyckas 14
22486 misslyckat 1
22487 misslyckats 9
22488 missnöjd 2
22489 missnöjda 1
22490 missnöje 4
22491 missriktade 1
22492 missta 1
22493 misstag 18
22494 misstagen 3
22495 misstaget 2
22496 misstankar 6
22497 misstanke 2
22498 misstar 3
22499 misstolkas 2
22500 misstro 5
22501 misstroende 1
22502 misstroendeförklaring 1
22503 misstroenderöst 1
22504 misstroendevotum 1
22505 misstrott 1
22506 misstänka 1
22507 misstänker 8
22508 misstänksamhet 3
22509 misstänksamt 1
22510 misstänkt 3
22511 misstänkta 1
22512 misstänkte 3
22513 missuppfattning 2
22514 missuppfattningar 2
22515 missöde 3
22516 missödet 1
22517 mist 3
22518 mista 1
22519 miste 7
22520 mister 1
22521 misär 1
22522 misären 2
22523 mitt 231
22524 mittemot 1
22525 mitten 6
22526 mittgången 1
22527 mittplatsen 1
22528 mix 4
22529 mixas 1
22530 mixtra 1
22531 mixtrade 1
22532 mjuk 4
22533 mjuka 3
22534 mjukade 1
22535 mjukades 1
22536 mjukare 1
22537 mjukat 1
22538 mjukhjärtad 1
22539 mjuklandning 1
22540 mjukt 3
22541 mjölk 1
22542 mjölke 1
22543 mjölkig 1
22544 mjölkprodukter 1
22545 mjölkpulver 2
22546 mobilisera 6
22547 mobiliserade 1
22548 mobiliserar 1
22549 mobiliseras 1
22550 mobiliserat 2
22551 mobiliserats 1
22552 mobilisering 3
22553 mobiliseringen 3
22554 mobilområdet 1
22555 mobiltelefoner 2
22556 mobiltelefonerna 1
22557 mobiltelefoni 1
22558 mobiltelefonin 1
22559 mod 8
22560 modebegreppet 1
22561 modell 27
22562 modellen 24
22563 modellens 1
22564 modeller 8
22565 modellerna 4
22566 modenyck 2
22567 modeordet 1
22568 moder 2
22569 moderat 1
22570 moderata 2
22571 modern 11
22572 moderna 21
22573 modernare 1
22574 modernisera 15
22575 moderniserade 1
22576 moderniseras 2
22577 modernisering 38
22578 moderniseringen 5
22579 moderniseringsprocess 2
22580 moderniseringsstrategi 1
22581 modernt 3
22582 moderskap 3
22583 modersmål 1
22584 modet 10
22585 modifiera 1
22586 modifierade 26
22587 modifierat 3
22588 modifierats 1
22589 modig 3
22590 modiga 8
22591 modige 2
22592 modigt 2
22593 modlösa 1
22594 mods 3
22595 modus 2
22596 mogen 3
22597 moget 1
22598 mogna 4
22599 mognad 2
22600 mognat 1
22601 moln 2
22602 molnen 3
22603 molnfria 1
22604 molnig 1
22605 moment 1
22606 momenten 1
22607 momspliktiga 1
22608 monetarism 3
22609 monetaristisk 1
22610 monetaristiska 1
22611 monetär 4
22612 monetära 17
22613 monitoring 1
22614 monokulturer 1
22615 monokulturerna 2
22616 monolog 1
22617 monopol 26
22618 monopolbildning 2
22619 monopolen 1
22620 monopolens 1
22621 monopolet 2
22622 monopolets 1
22623 monopolfrågor 1
22624 monopolföretag 1
22625 monopolföretags 1
22626 monopolintressen 1
22627 monopoliserade 3
22628 monopoliserats 1
22629 monopoliska 1
22630 monopolmarknader 1
22631 monopolrättigheter 1
22632 monopolsituation 1
22633 monopolställning 1
22634 monster 1
22635 monsterhustrun 1
22636 monstermannen 1
22637 monstermasken 1
22638 monsterälskarinnan 1
22639 monterat 1
22640 mopp 1
22641 moppen 1
22642 mor 33
22643 moral 5
22644 moralen 3
22645 moralisk 2
22646 moraliska 7
22647 moraliskt 4
22648 moralism 1
22649 moratorium 1
22650 morbror 17
22651 morbrors 1
22652 mord 10
22653 mordbränder 1
22654 morden 1
22655 mordet 2
22656 mordförsöken 1
22657 mordiska 1
22658 morgnar 2
22659 morgon 127
22660 morgon- 1
22661 morgondagen 2
22662 morgondagens 7
22663 morgonen 8
22664 morgonregn 1
22665 morgons 1
22666 morgonsolen 1
22667 morgonteet 1
22668 morgontimmen 1
22669 mormodern 1
22670 mormonmissionär 1
22671 mormor 6
22672 morot 1
22673 morrade 1
22674 morron 1
22675 morronen 1
22676 mors 3
22677 morse 22
22678 moskiter 1
22679 moskéns 1
22680 moster 8
22681 mot 769
22682 motarbeta 6
22683 motarbetar 1
22684 motbjudande 2
22685 motgångar 1
22686 motgångarna 1
22687 motion 2
22688 motionen 1
22689 motioner 2
22690 motiv 9
22691 motivation 4
22692 motivationen 2
22693 motiven 3
22694 motivera 8
22695 motiverad 2
22696 motiverade 5
22697 motiverades 1
22698 motiverar 9
22699 motiveras 2
22700 motiverat 1
22701 motiverats 1
22702 motivering 7
22703 motiveringar 2
22704 motiveringen 5
22705 motivet 2
22706 motljus 2
22707 motor 3
22708 motorcyklar 3
22709 motorcyklarna 1
22710 motorer 1
22711 motorerna 3
22712 motorindustrin 2
22713 motorister 1
22714 motorn 3
22715 motorns 2
22716 motorväg 2
22717 motorvägar 1
22718 motpart 2
22719 motparten 2
22720 motpartens 1
22721 motparter 1
22722 motpartsmedel 1
22723 motsats 24
22724 motsatsen 11
22725 motsatser 1
22726 motsatsförhållande 1
22727 motsatsställning 1
22728 motsatt 9
22729 motsatta 12
22730 motsatte 3
22731 motstridig 1
22732 motstridiga 8
22733 motstridigheter 2
22734 motsträvig 1
22735 motsträvigt 1
22736 motstycke 6
22737 motstånd 10
22738 motståndare 13
22739 motståndarna 1
22740 motståndet 5
22741 motståndsrörelser 1
22742 motstår 2
22743 motsvara 2
22744 motsvarade 1
22745 motsvarades 1
22746 motsvarande 31
22747 motsvarar 22
22748 motsvaras 1
22749 motsvarats 1
22750 motsvarighet 5
22751 motsvarigheter 2
22752 motsäga 1
22753 motsägande 2
22754 motsägas 1
22755 motsägelse 7
22756 motsägelsefull 1
22757 motsägelsefulla 7
22758 motsägelsefullt 8
22759 motsägelsens 1
22760 motsägelser 3
22761 motsägelserna 1
22762 motsätta 3
22763 motsätter 17
22764 motsättning 8
22765 motsättningar 16
22766 motsättningarna 5
22767 motsättningen 1
22768 motta 1
22769 mottaga 1
22770 mottagande 6
22771 mottagandet 4
22772 mottagare 1
22773 mottagarlandet 2
22774 mottagarlandets 2
22775 mottagarländerna 2
22776 mottagarländernas 1
22777 mottagarna 2
22778 mottagarområden 1
22779 mottagarområdena 1
22780 mottagarprogrammet 1
22781 mottagit 11
22782 mottagits 4
22783 mottagna 1
22784 mottagning 1
22785 mottagningar 1
22786 mottagningarna 1
22787 mottagningsanläggning 1
22788 mottagningsanläggningar 3
22789 mottagningsanläggningen 1
22790 mottagningsanordningar 7
22791 mottagningsanordningarna 1
22792 mottagningsbevis 1
22793 mottagningsceremoni 1
22794 mottagningsförhållanden 1
22795 mottar 1
22796 motto 1
22797 mottog 3
22798 mottogs 2
22799 motverka 9
22800 motverkar 2
22801 motvikt 2
22802 motvilja 1
22803 motvilligt 3
22804 motvärn 1
22805 motåtgärd 1
22806 motåtgärder 5
22807 moçambikier 2
22808 moçambikierna 1
22809 moçambikiska 3
22810 mr 23
22811 mrs 14
22812 muddermassorna 1
22813 muddras 1
22814 mugglare 2
22815 mugglarkvinna 1
22816 mugglarpengar 1
22817 mugglarägare 1
22818 mullrande 1
22819 mullvad 1
22820 multi-etniska 1
22821 multi-etniskt 1
22822 multietnisk 1
22823 multietniska 3
22824 multietniskt 2
22825 multilateral 2
22826 multilaterala 7
22827 multinationell 1
22828 multinationella 16
22829 multinationellt 1
22830 multipliceras 1
22831 multiplikatoreffekt 2
22832 multiplikatoreffekten 1
22833 mumifierade 1
22834 mumla 1
22835 mumlade 4
22836 mumlande 1
22837 mun 9
22838 munnen 5
22839 muntera 1
22840 munterhet 1
22841 muntert 1
22842 muntlig 2
22843 muntliga 23
22844 muntligen 1
22845 muntligt 4
22846 muntra 1
22847 mur 3
22848 murad 1
22849 murar 3
22850 muren 1
22851 museifartyg 1
22852 museifartygen 1
22853 muselmansk 1
22854 museum 1
22855 musik 6
22856 musikanter 1
22857 musiken 3
22858 musiker 1
22859 muskler 1
22860 muskulös 1
22861 muslim 1
22862 mussel- 3
22863 musselodlare 2
22864 must 1
22865 mustasch 1
22866 mustascher 1
22867 mustascherna 1
22868 muta 1
22869 mutgle-baiting 1
22870 mutor 1
22871 muttrade 3
22872 muttrande 2
22873 mycken 3
22874 mycket 1417
22875 mygg 1
22876 myggen 1
22877 myggor 1
22878 myllan 1
22879 myllrade 2
22880 myllrande 1
22881 myllrar 1
22882 myndiga 1
22883 myndigförklarade 1
22884 myndighet 27
22885 myndigheten 30
22886 myndighetens 16
22887 myndigheter 68
22888 myndigheterna 105
22889 myndigheternas 13
22890 myndigheters 4
22891 myndighetsförfaranden 1
22892 myndighetskrångel 1
22893 myndighetsåtgärder 1
22894 mynna 4
22895 mynning 2
22896 mynningarna 1
22897 mynningen 3
22898 mynningsområde 1
22899 mynningsområdet 1
22900 mynt 4
22901 mynten 2
22902 myror 4
22903 mysteriejakt 1
22904 mysterier 1
22905 mysterium 5
22906 mystiska 2
22907 mytiskt 1
22908 mäkleriverksamhet 1
22909 mäkta 1
22910 mäktig 1
22911 mäktiga 2
22912 mäktigaste 1
22913 män 85
22914 mängd 34
22915 mängden 7
22916 mängder 12
22917 mängdfunktionerna 1
22918 mängdfunktionsreferens 1
22919 männen 22
22920 männens 3
22921 människa 14
22922 människan 14
22923 människans 9
22924 människo- 1
22925 människoben 1
22926 människoföda 2
22927 människoföraktande 1
22928 människoförföljande 1
22929 människohandel 3
22930 människoknotor 1
22931 människokompost 1
22932 människokännedom 1
22933 människokärlek 1
22934 människoliv 10
22935 människomassan 1
22936 människomyller 1
22937 människonaglar 1
22938 människor 234
22939 människorna 51
22940 människornas 5
22941 människors 35
22942 människorätten 1
22943 människorättskommissionerna 1
22944 människorättsnarcissismen 1
22945 människorättsnivån 1
22946 människorättsorganisationer 2
22947 människorättspolitik 5
22948 människorättspolitiken 3
22949 människosläktet 2
22950 människosmugglarnas 1
22951 människosmuggling 1
22952 människosyn 1
22953 människovänlig 1
22954 människovärdet 1
22955 människovärdiga 2
22956 människovärdigt 1
22957 mäns 2
22958 mänsklig 15
22959 mänskliga 247
22960 mänskligheten 6
22961 mänskligt 6
22962 märk 1
22963 märka 6
22964 märkas 1
22965 märkbar 5
22966 märkbara 3
22967 märkbart 2
22968 märke 19
22969 märken 5
22970 märker 4
22971 märkesgrupperna 1
22972 märklig 4
22973 märkliga 4
22974 märkligare 1
22975 märkligheter 1
22976 märkligt 6
22977 märkning 13
22978 märkningen 4
22979 märks 1
22980 märkt 2
22981 märkte 3
22982 märkvärdig 1
22983 märkvärdiga 1
22984 märkvärdigt 4
22985 mäss 1
22986 mässan 1
22987 mässing-tråd 1
22988 mässingsinstrument 1
22989 mästerverk 4
22990 mäta 9
22991 mätare 3
22992 mätas 5
22993 mätbara 2
22994 mäter 1
22995 mätningar 1
22996 mäts 3
22997 mätt 2
22998 mätte 1
22999 mättes 1
23000 må 17
23001 måfå 1
23002 måhända 7
23003 mål 283
23004 mål-2-området 1
23005 måla 3
23006 målade 3
23007 målar 1
23008 målarfärg 1
23009 målas 1
23010 målat 1
23011 målats 2
23012 målen 48
23013 målens 1
23014 målet 62
23015 målformat 1
23016 målgrupp 2
23017 målgrupper 1
23018 målgången 1
23019 målinriktad 1
23020 målinriktade 2
23021 målinriktat 5
23022 mållösa 1
23023 målmedvetet 3
23024 målområdena 1
23025 målområdet 1
23026 målsättning 25
23027 målsättningar 25
23028 målsättningarna 16
23029 målsättningen 16
23030 måltid 3
23031 måltidens 1
23032 mån 31
23033 mån. 1
23034 måna 3
23035 månad 33
23036 månaden 17
23037 månader 92
23038 månaderna 35
23039 månaders 1
23040 månads 2
23041 månadslånga 1
23042 månadsvisa 1
23043 månatliga 1
23044 månbelyst 1
23045 måndag 7
23046 måndagar 1
23047 måndagen 2
23048 måndags 11
23049 månde 1
23050 måne 1
23051 många 577
23052 mångbesjungna 1
23053 mångfald 25
23054 mångfalden 16
23055 mångfaldig 1
23056 mångfaldiga 4
23057 mångfaldigandet 1
23058 mångfaldigas 1
23059 mångfaldigt 2
23060 mångformiga 1
23061 mångfunktionell 1
23062 mångfärgad 1
23063 mångkulturella 2
23064 mångkunnig 1
23065 mångnationellt 1
23066 mångsidighet 1
23067 mångsidigt 4
23068 mångskiftande 1
23069 mångt 2
23070 mångtaliga 1
23071 mångtydiga 1
23072 mångåriga 2
23073 månljuset 1
23074 månsken 1
23075 mår 3
23076 måste 1985
23077 mått 9
23078 måtte 2
23079 måttenhet 2
23080 måttet 1
23081 måttfulla 1
23082 måttfullhet 1
23083 måttlig 1
23084 måtto 7
23085 måttstock 4
23086 måttstocken 1
23087 möblemanget 1
23088 möbler 4
23089 möblerad 1
23090 möblerna 1
23091 möda 5
23092 mödan 1
23093 mödosam 1
23094 mödosamma 1
23095 mödosamt 1
23096 mödrar 2
23097 möjlig 15
23098 möjliga 63
23099 möjligen 12
23100 möjliggjorde 1
23101 möjliggjort 3
23102 möjliggör 13
23103 möjliggöra 23
23104 möjliggörs 2
23105 möjlighet 130
23106 möjligheten 55
23107 möjligheter 129
23108 möjligheterna 22
23109 möjligheternas 4
23110 möjligheteten 1
23111 möjligt 340
23112 möjligtvis 3
23113 mönster 4
23114 mönsterbild 1
23115 mönsterskydd 1
23116 mönstring 1
23117 mördade 1
23118 mördades 2
23119 mördande 2
23120 mördar 1
23121 mördare 2
23122 mördaren 2
23123 mördas 1
23124 mördat 2
23125 mördats 2
23126 mörk 4
23127 mörka 18
23128 mörkare 2
23129 mörkblond 1
23130 mörkblå 1
23131 mörker 4
23132 mörkgröna 1
23133 mörklägga 1
23134 mörknade 1
23135 mörkret 14
23136 mörkrets 2
23137 mörkrött 1
23138 mörkt 7
23139 möta 29
23140 mötas 1
23141 möte 48
23142 möten 14
23143 mötena 2
23144 möter 7
23145 mötes 6
23146 mötespunkt 1
23147 mötet 22
23148 möts 3
23149 mött 1
23150 mötte 2
23151 möttes 3
23152 mötts 2
23153 müssen 2
23154 n 3
23155 nackdel 8
23156 nackdelar 7
23157 nacke 1
23158 nacken 4
23159 nagel 1
23160 naglar 1
23161 naiva 1
23162 naivitet 1
23163 naivt 1
23164 nakna 2
23165 nallebjörn 1
23166 namn 52
23167 namnen 1
23168 namnet 26
23169 namnfrågan 1
23170 namnlös 1
23171 namnlösa 1
23172 namnteckning 2
23173 namnupprop 6
23174 nappat 1
23175 narkotika 3
23176 narkotikabekämpning 1
23177 narkotikahandel 1
23178 narkotikahandeln 1
23179 narkotikamissbrukare 1
23180 narkotikan 1
23181 narkotikaproblematiken 1
23182 narkotikasmuggling 2
23183 narrarnas 1
23184 nation 5
23185 national 1
23186 national-socialistiska 1
23187 nationalekonomin 1
23188 nationalekonomisk 1
23189 nationalekonomiska 3
23190 nationalekonomiskt 2
23191 nationalförsamling 1
23192 nationalförsamlingen 3
23193 nationaliseringsprocess 1
23194 nationalism 4
23195 nationalismens 1
23196 nationalister 1
23197 nationalisterna 1
23198 nationalistiska 1
23199 nationalitet 5
23200 nationaliteter 3
23201 nationalklänning 1
23202 nationalliberaler 1
23203 nationalräkenskapssystemet 6
23204 nationalsocialismen 1
23205 nationalstaten 2
23206 nationalstatens 1
23207 nationalstater 2
23208 nationalstaterna 1
23209 nationalsången 1
23210 nationell 46
23211 nationella 260
23212 nationellt 13
23213 nationen 1
23214 nationens 2
23215 nationer 12
23216 nationerna 25
23217 nationernas 39
23218 nationsgränser 2
23219 nationsregionerna 1
23220 nationsskapande 1
23221 nationsspecifika 1
23222 natt 5
23223 nattblommor 1
23224 natten 20
23225 nattens 2
23226 nattetid 1
23227 nattfjärilar 1
23228 nattfjärilsmjuka 1
23229 nattliga 2
23230 nattlinne 1
23231 nattsaga 1
23232 nattsammanträden 1
23233 nattsammanträdenas 1
23234 nattsäck 1
23235 nattupplagan 1
23236 nattvagabonderande 1
23237 nattvinden 1
23238 nattväskan 1
23239 natur 29
23240 natur- 3
23241 natura 1
23242 naturarvet 1
23243 naturen 19
23244 naturens 2
23245 naturfenomen 1
23246 naturkatastrof 2
23247 naturkatastrofen 2
23248 naturkatastrofer 17
23249 naturlig 8
23250 naturliga 19
23251 naturligt 16
23252 naturligtvis 237
23253 naturnätverket 1
23254 naturnödvändighet 1
23255 naturområden 2
23256 naturresurs 3
23257 naturresurser 4
23258 naturresurserna 5
23259 naturskydd 1
23260 naturskyddspolitiken 1
23261 naturtillgångar 4
23262 naturvetenskaplig 1
23263 naturvidrigt 1
23264 navajoindianerna 1
23265 navajoreservatet 1
23266 navigationssektionen 1
23267 navigerat 1
23268 nazism 2
23269 nazismen 4
23270 nazismens 1
23271 nazist 3
23272 nazistflirtande 1
23273 nazistisk 1
23274 ne 1
23275 necessär 2
23276 necessären 1
23277 ned 65
23278 nedan 1
23279 nedanför 5
23280 nedbrytningen 1
23281 nedbrända 1
23282 nedbäddad 1
23283 neddragna 1
23284 neddragningar 1
23285 nederbörd 1
23286 nederbörden 2
23287 nederlag 2
23288 nederländare 1
23289 nederländsk 11
23290 nederländsk-brittisk-skandinavisk 1
23291 nederländska 15
23292 nedersta 1
23293 nedför 1
23294 nedgång 3
23295 nedgången 2
23296 nedifrån 1
23297 nedkomma 1
23298 nedkomst 1
23299 nedlagd 1
23300 nedlagda 1
23301 nedläggning 2
23302 nedläggningar 2
23303 nedläggningen 1
23304 nedlåta 1
23305 nedlåtande 1
23306 nedmontera 1
23307 nedmontering 2
23308 nedmonterings- 1
23309 nedre 1
23310 nedrullningsbara 1
23311 nedrustning 1
23312 nedrustningen 1
23313 nedskräpningsproblem 1
23314 nedskärning 2
23315 nedskärningar 6
23316 nedskärningspolitik 1
23317 nedsmutsade 2
23318 nedsmutsning 3
23319 nedsmutsningen 4
23320 nedströms 5
23321 nedstämd 1
23322 nedstängning 1
23323 nedstängningsplaner 1
23324 nedsänkt 1
23325 nedsättande 1
23326 nedtecknat 1
23327 nedvärdera 1
23328 nedvärderas 1
23329 nedåt 6
23330 negativ 14
23331 negativa 38
23332 negativism 1
23333 negativt 21
23334 neger 1
23335 negligera 1
23336 nej 26
23337 nejlikor 1
23338 neka 3
23339 nekad 1
23340 nekande 1
23341 nekas 5
23342 neo-liberalism 1
23343 neofascistiska 2
23344 neoklassiska 1
23345 neokolonial 1
23346 neokolonialismen 1
23347 neokolonialistiska 1
23348 neonazistiskt 1
23349 neonlampor 1
23350 nepotism 5
23351 ner 97
23352 nerdrogad 1
23353 nere 17
23354 nerför 12
23355 nerhukade 1
23356 nerver 1
23357 nervkrig 1
23358 nervpåfrestande 1
23359 nervös 3
23360 nervösa 1
23361 nervöst 3
23362 netto 1
23363 nettoupplåning 1
23364 nettoökning 1
23365 neutral 1
23366 neutrala 2
23367 neutraliserar 1
23368 neutraliseras 1
23369 neutralitet 1
23370 neutralt 2
23371 neutre 2
23372 new 6
23373 ni 833
23374 nickade 4
23375 nigerianska 1
23376 niggrer 1
23377 nihilo-rätt 1
23378 nikotinproblemen 1
23379 nimbus 1
23380 nio 18
23381 nionde 2
23382 nioåring 1
23383 nischer 1
23384 nit 1
23385 nitratdirektivet 1
23386 nittiotalet 1
23387 nitton 2
23388 nittonhundra 1
23389 nittonhundrafyrtitalet 1
23390 nittonhundratalet 1
23391 nittonhundratalets 1
23392 nivå 169
23393 nivåer 23
23394 nivåerna 2
23395 nivån 15
23396 njuta 2
23397 njuter 2
23398 njutning 3
23399 njöt 4
23400 nn 1
23401 no 6
23402 nobelpristagaren 1
23403 nog 56
23404 noga 37
23405 noggrann 7
23406 noggranna 5
23407 noggrannare 4
23408 noggrannhet 4
23409 noggrannheten 1
23410 noggrant 29
23411 noll 17
23412 noll-alternativet 1
23413 nollgradig 3
23414 nollgränsvärde 1
23415 nollkravet 1
23416 nollning 1
23417 nollnivå 1
23418 nollnivårisk 1
23419 nollor 1
23420 nollrisk 1
23421 nollstrecket 1
23422 nollställda 1
23423 nollutsläpp 2
23424 nollårig 1
23425 nominell 2
23426 nominella 2
23427 nominera 4
23428 nominerade 1
23429 nominerar 1
23430 nomineras 1
23431 nomineringen 1
23432 non 4
23433 nonchalansen 1
23434 nonchalant 1
23435 nonchalerade 2
23436 nonsens 2
23437 nonsensord 1
23438 nord 1
23439 nord-syd 2
23440 nordafrikanska 3
23441 nordamerikanerna 1
23442 nordamerikanska 6
23443 nordeuropeiska 1
23444 nordirländare 1
23445 nordirländska 1
23446 nordisk 1
23447 nordiska 4
23448 nordkusten 1
23449 nordlig 1
23450 nordliga 6
23451 nordtyska 1
23452 nordvästra 4
23453 norm 2
23454 normal 6
23455 normala 10
23456 normaliserades 1
23457 normalisering 5
23458 normaliseringen 2
23459 normalitet 1
23460 normalt 17
23461 normativ 1
23462 normativt 2
23463 normen 1
23464 normer 36
23465 normerna 15
23466 normgivande 1
23467 norr 9
23468 norr-söder 1
23469 norra 25
23470 norrmännens 1
23471 norrut 2
23472 norska 2
23473 norskt 1
23474 nos 1
23475 noshörning 1
23476 nosspetsen 1
23477 nostrum 1
23478 not 3
23479 notan 1
23480 notera 23
23481 noterade 6
23482 noterades 1
23483 noterar 28
23484 noteras 3
23485 noterat 17
23486 noterna 1
23487 notis 1
23488 november 30
23489 nr 81
23490 nu 713
23491 nuet 2
23492 nuets 1
23493 null-värden 5
23494 nulla 1
23495 nullitetssanktionen 1
23496 nullvärde 1
23497 nuläget 5
23498 numer 1
23499 numera 19
23500 numerära 1
23501 nummer 12
23502 numreringen 1
23503 numret 6
23504 nunnor 1
23505 nutida 1
23506 nuvarande 145
23507 ny 174
23508 nya 630
23509 nyanlända 1
23510 nyans 1
23511 nyansera 1
23512 nyanserad 1
23513 nyanserna 1
23514 nyanställda 2
23515 nyanställningar 1
23516 nyare 1
23517 nyaste 1
23518 nybildande 1
23519 nybilsköparna 1
23520 nybilspriset 1
23521 nybyggarens 1
23522 nybyggets 1
23523 nyckel 2
23524 nyckelfaktor 1
23525 nyckelfråga 3
23526 nyckelfrågan 1
23527 nyckelfrågor 1
23528 nyckelfrågorna 1
23529 nyckelfunktioners 1
23530 nyckeln 6
23531 nyckelområden 1
23532 nyckelord 1
23533 nyckelorden 1
23534 nyckelordet 1
23535 nyckelproblem 2
23536 nyckelpunkter 1
23537 nyckelroll 3
23538 nyckelsektor 1
23539 nyckelåtgärder 1
23540 nycklar 1
23541 nycklarna 1
23542 nydanande 6
23543 nye 3
23544 nyetableringar 1
23545 nyexaminerad 1
23546 nyfascister 1
23547 nyfattigdom 1
23548 nyfiken 4
23549 nyfiket 1
23550 nyfikna 1
23551 nyföretagarvänlig 1
23552 nyförvärvade 1
23553 nygift 1
23554 nyhet 6
23555 nyheten 1
23556 nyheter 15
23557 nyheterna 9
23558 nyhetsinslag 1
23559 nyhetsprogrammet 1
23560 nyhetsrapporterna 1
23561 nykomlingar 1
23562 nykomlingarna 1
23563 nyktert 3
23564 nyktra 1
23565 nylansera 1
23566 nylansering 1
23567 nylanseringen 1
23568 nyliberal 2
23569 nyliberala 2
23570 nyliberalt 1
23571 nyligen 87
23572 nylon 1
23573 nylonet 1
23574 nylonspetsar 1
23575 nylontrosornas 1
23576 nynazism 1
23577 nynazismen 1
23578 nynazist 1
23579 nynazister 2
23580 nynazistiska 1
23581 nypa 1
23582 nypan 1
23583 nyplanteringen 1
23584 nyskapande 3
23585 nyss 46
23586 nystart 1
23587 nytt 155
23588 nytta 55
23589 nyttan 5
23590 nyttig 7
23591 nyttiga 8
23592 nyttighet 1
23593 nyttigt 4
23594 nyttjande 1
23595 nyttoanalys 1
23596 nyttobruk 1
23597 nyttofordon 9
23598 nytänkande 3
23599 nyval 1
23600 nyvald 1
23601 nyvalda 1
23602 nyvalde 1
23603 nyårsaftonen 1
23604 näbbig 1
23605 nämligen 204
23606 nämna 63
23607 nämnare 1
23608 nämnaren 2
23609 nämnas 3
23610 nämnda 17
23611 nämnde 45
23612 nämndes 9
23613 nämner 25
23614 nämns 24
23615 nämnt 27
23616 nämnts 20
23617 nämnvärd 1
23618 nämnvärda 1
23619 nämnvärt 1
23620 när 1122
23621 nära 83
23622 närapå 1
23623 närbelägna 2
23624 närbesläktad 1
23625 närbesläktade 1
23626 närekonomi 1
23627 närhelst 1
23628 närhet 1
23629 närheten 16
23630 närhetsamtal 1
23631 näring 1
23632 näringar 3
23633 näringsgren 3
23634 näringsgrenen 1
23635 näringsidkare 1
23636 näringskedja 1
23637 näringskedjan 1
23638 näringsliv 1
23639 näringslivet 14
23640 näringslivets 5
23641 näringslivsaktörer 1
23642 näringsrik 1
23643 näringsstrukturen 1
23644 näringstillskott 1
23645 näringsvärden 1
23646 närliggande 1
23647 närma 10
23648 närmade 3
23649 närmande 10
23650 närmanden 1
23651 närmandet 1
23652 närmar 8
23653 närmare 51
23654 närmast 16
23655 närmaste 53
23656 närmsta 1
23657 närområdet 2
23658 närpolisen 1
23659 närpoliser 1
23660 närpolissystem 1
23661 närstående 4
23662 närsynt 2
23663 närvara 6
23664 närvarade 1
23665 närvarande 127
23666 närvarar 1
23667 närvaro 26
23668 närvaron 6
23669 näsa 5
23670 näsan 8
23671 näsborrar 1
23672 näsdukar 1
23673 näsduken 1
23674 näst 1
23675 nästa 98
23676 nästan 97
23677 nästkommande 1
23678 näsvingarna 1
23679 nät 12
23680 näten 5
23681 nätens 1
23682 nätet 3
23683 nätstrukturer 1
23684 nätt 2
23685 nätter 3
23686 nätterna 1
23687 nätverk 13
23688 nätverken 3
23689 nätverkens 2
23690 nätverket 2
23691 nätverkslicens 1
23692 nätverkslicensavtal 1
23693 nätverkslicensen 1
23694 nätverkssamhället 1
23695 nå 70
23696 nåbar 2
23697 nåd 2
23698 nådde 6
23699 nåddes 2
23700 nåden 1
23701 någon 468
23702 någons 1
23703 någonsin 33
23704 någonstans 30
23705 någonting 112
23706 någonvart 1
23707 någorlunda 2
23708 något 638
23709 någotdera 1
23710 några 464
23711 nåja 1
23712 nål 1
23713 nån 4
23714 nånsin 3
23715 nånstans 4
23716 nånting 3
23717 når 9
23718 nås 4
23719 nåt 7
23720 nått 23
23721 nåtts 1
23722 nöd 3
23723 nödbedd 1
23724 nöden 2
23725 nödens 1
23726 nödfall 1
23727 nödgas 2
23728 nödhjälp 4
23729 nödhjälpen 1
23730 nödinsatser 1
23731 nödlösning 1
23732 nödraketer 1
23733 nödreparationer 1
23734 nödsituation 2
23735 nödsituationen 1
23736 nödsituationer 1
23737 nödsituationsfasen 1
23738 nödställda 1
23739 nödtorftiga 1
23740 nödvändig 51
23741 nödvändiga 85
23742 nödvändigare 1
23743 nödvändiggör 1
23744 nödvändighet 12
23745 nödvändigheten 18
23746 nödvändigheterna 1
23747 nödvändighetsperspektiv 1
23748 nödvändigt 205
23749 nödvändigtvis 19
23750 nödåtgärder 1
23751 nöja 20
23752 nöjaktig 1
23753 nöjaktigt 1
23754 nöjd 14
23755 nöjda 16
23756 nöjde 1
23757 nöje 14
23758 nöjer 6
23759 nöjesbåtar 1
23760 nöjessökande 1
23761 nöjet 7
23762 nöjsam 1
23763 nöjt 2
23764 nöt 1
23765 nötkreatur 1
23766 nötkött 7
23767 nötkötts- 1
23768 nötköttsöverskott 1
23769 nötskal 2
23770 nött 1
23771 nötter 1
23772 nötterna 1
23773 nöttköttslager 1
23774 o 3
23775 o.s.v. 2
23776 oacceptabel 19
23777 oacceptabelt 31
23778 oacceptabla 17
23779 oaktat 2
23780 oanmälda 3
23781 oansenligt 1
23782 oanständiga 1
23783 oansvariga 3
23784 oansvarighet 6
23785 oansvarigheten 1
23786 oanvända 1
23787 oanvändbar 2
23788 oanvändbart 1
23789 oartig 1
23790 oavbruten 2
23791 oavbrutet 2
23792 oavbrutna 1
23793 oavhängighet 2
23794 oavhängighetsförklaringen 2
23795 oavsett 42
23796 oavsiktlig 1
23797 oavsiktliga 3
23798 oavsiktligt 1
23799 oavslutade 1
23800 oavvislig 1
23801 obalans 6
23802 obalansen 5
23803 obalanser 2
23804 obalanserna 2
23805 obarmhärtiga 1
23806 obarmhärtigt 1
23807 obeboelig 1
23808 obefintliga 2
23809 obefläckad 2
23810 obefogat 2
23811 obegriplig 2
23812 obegripliga 1
23813 obegripligt 3
23814 obegränsad 6
23815 obegränsat 1
23816 obehag 1
23817 obehagliga 2
23818 obehagligt 4
23819 obekant 2
23820 obekanta 1
23821 obekväm 1
23822 obekväma 1
23823 obekymrad 1
23824 obekymrade 2
23825 obemannad 1
23826 obemärkt 3
23827 obemärkthet 1
23828 oberoende 85
23829 oberoendes 1
23830 oberoendet 1
23831 oberättigad 1
23832 oberättigat 1
23833 oberörd 2
23834 oberörda 1
23835 obestridlig 1
23836 obestridliga 2
23837 obestämd 4
23838 obesvarad 1
23839 obesvarade 3
23840 obesvarbara 1
23841 obesvärade 1
23842 obetalda 2
23843 obetydlig 2
23844 obetydligt 1
23845 obevakade 1
23846 obevekliga 1
23847 obeveklighet 1
23848 obeväpnade 1
23849 obildad 1
23850 objekt 11
23851 objektbibliotek 1
23852 objektdefinitioner 1
23853 objekten 1
23854 objektet 2
23855 objektets 1
23856 objektiv 3
23857 objektiva 5
23858 objektivt 7
23859 oblandad 1
23860 obligationer 1
23861 obligationsmarknaderna 1
23862 obligatorisk 13
23863 obligatoriska 12
23864 obligatoriskt 4
23865 obligatorium 1
23866 obrukbart 1
23867 observation 2
23868 observationerna 1
23869 observatorium 1
23870 observatory 2
23871 observatörens 1
23872 observatörer 6
23873 observatörerna 1
23874 observera 2
23875 observerats 1
23876 obsolet 1
23877 obundna 3
23878 obönhörligt 1
23879 oceanen 1
23880 oceanerna 2
23881 oceanernas 1
23882 och 15689
23883 också 1597
23884 ockupanten 1
23885 ockupation 2
23886 ockupationen 4
23887 ockupationsmakt 1
23888 ockupationsstyrkorna 1
23889 ockuperade 15
23890 ockuperades 1
23891 ockuperande 1
23892 ockuperas 1
23893 ockuperat 1
23894 odds 1
23895 odefinierade 1
23896 odefinierbart 1
23897 odelad 1
23898 odelade 1
23899 odelbara 1
23900 odemokratiska 2
23901 odifferentierad 1
23902 odiskutabel 1
23903 odiskutabelt 1
23904 odjur 2
23905 odla 4
23906 odlad 1
23907 odlar 1
23908 odlare 1
23909 odlarna 3
23910 odling 3
23911 odlingar 7
23912 odlingarna 1
23913 odlingen 1
23914 odlingsmarker 1
23915 odlingsplatser 1
23916 odugliga 1
23917 odödliga 1
23918 oeftergivligt 1
23919 oegennyttiga 2
23920 oegentlig 1
23921 oegentliga 1
23922 oegentlighet 2
23923 oegentligheter 3
23924 oegentligheterna 1
23925 oegentligt 1
23926 oekonomisk 1
23927 oekonomiskt 1
23928 oemotståndlig 1
23929 oemotståndligt 1
23930 oemotsägligt 1
23931 oenighet 5
23932 oenigheten 1
23933 oenigheterna 1
23934 oense 5
23935 oerhörd 4
23936 oerhörda 5
23937 oerhört 25
23938 oersättliga 1
23939 oetiska 1
23940 of 14
23941 ofantlig 1
23942 ofantliga 5
23943 ofantligt 1
23944 ofarlig 3
23945 ofarligt 1
23946 ofattbara 3
23947 ofattbart 1
23948 ofelbara 1
23949 offensiv 2
23950 offensiva 1
23951 offensiven 1
23952 offensivt 3
23953 offentlig 38
23954 offentliga 152
23955 offentligen 1
23956 offentliggjorda 1
23957 offentliggjorde 5
23958 offentliggjordes 2
23959 offentliggjort 3
23960 offentliggjorts 4
23961 offentliggör 2
23962 offentliggöra 7
23963 offentliggörande 1
23964 offentliggörandet 2
23965 offentliggöras 6
23966 offentliggörs 5
23967 offentlighet 2
23968 offentligheten 2
23969 offentlighetens 2
23970 offentlighetsförordningen 1
23971 offentlighetskampanj 1
23972 offentlighetsprincip 1
23973 offentligpolitiska 1
23974 offentligt 16
23975 offer 32
23976 officerare 1
23977 officiell 1
23978 officiella 20
23979 officiellt 7
23980 offra 1
23981 offrade 1
23982 offrades 1
23983 offrar 1
23984 offras 4
23985 offren 25
23986 offrens 4
23987 offret 2
23988 oflexibilitet 1
23989 oformaterad 1
23990 oframkomlig 1
23991 ofred 1
23992 ofruktbart 1
23993 ofruktsamhet 1
23994 ofrånkomligen 3
23995 ofrånkomligt 3
23996 ofta 160
23997 oftare 14
23998 oftast 7
23999 ofullkomlighet 1
24000 ofullkomligt 1
24001 ofullständig 3
24002 ofullständiga 4
24003 ofullständigt 1
24004 ofärdig 1
24005 oförblommerat 1
24006 ofördelaktiga 1
24007 ofördelaktigaste 1
24008 ofördelaktigt 2
24009 oförenlig 2
24010 oförenliga 2
24011 oförenlighet 1
24012 oförenligt 4
24013 oförklarat 1
24014 oförklarlig 2
24015 oförklarliga 1
24016 oförklarligt 1
24017 oförlåtlig 1
24018 oförlåtligt 2
24019 oförmåga 7
24020 oförmågan 3
24021 oförmögen 3
24022 oförmögna 1
24023 oförnekligen 1
24024 oförnuftigt 1
24025 oförorenade 1
24026 oförsiktigt 2
24027 oförskämda 1
24028 oförståeligt 2
24029 oförsvarlig 2
24030 oförsvarligt 1
24031 oförtjänt 1
24032 oförtrutet 1
24033 oförtröttat 1
24034 oförutsägbar 1
24035 oföränderlig 3
24036 oföränderliga 1
24037 oföränderlighet 1
24038 oförändrad 2
24039 oförändrade 4
24040 oförändrat 1
24041 ogenomförbar 2
24042 ogenomskinligheten 1
24043 ogenomträngligt 1
24044 ogifta 1
24045 ogillande 1
24046 ogiltigförklarades 1
24047 ogrundad 1
24048 ogrundat 1
24049 ogräs 2
24050 ogynnsam 1
24051 ogynnsamma 2
24052 ogynnsamt 1
24053 ohejdad 1
24054 ohjälpligt 2
24055 ohyggliga 1
24056 ohyggligt 1
24057 ohygienisk 2
24058 ohyra 1
24059 ohälsa 1
24060 ohälsosamma 2
24061 ohälsosamt 1
24062 ohämmad 2
24063 ohämmade 3
24064 ohållbar 1
24065 ohållbara 1
24066 ohållbart 1
24067 ohörsamma 1
24068 ohövlig 2
24069 ohövliga 1
24070 oidily 1
24071 oigenkännelighet 1
24072 oinskränkt 1
24073 oinskränkta 2
24074 oinspelade 1
24075 ointelligent 1
24076 ointressant 1
24077 ointresse 3
24078 ointresserad 1
24079 ointresset 1
24080 ojordiska 1
24081 ojämförbar 1
24082 ojämlik 1
24083 ojämlikhet 9
24084 ojämlikheten 3
24085 ojämlikheter 3
24086 ojämlikheterna 1
24087 ojämn 2
24088 ojämna 2
24089 ojämnt 3
24090 okaraktäristiskt 1
24091 oket 1
24092 oklanderlig 2
24093 oklanderliga 1
24094 oklanderligt 1
24095 oklar 4
24096 oklara 4
24097 oklarhet 4
24098 oklarheter 5
24099 oklart 5
24100 oklok 1
24101 oklokt 1
24102 okomplicerad 1
24103 okomplicerade 2
24104 okongena 1
24105 okonstlad 1
24106 okontrollerad 4
24107 okontrollerade 3
24108 okontrollerat 1
24109 okontrollerbar 1
24110 okontrollerbara 1
24111 okritiska 1
24112 okritiskt 3
24113 okränkbara 2
24114 okränkbarheten 1
24115 oktaverna 1
24116 oktober 24
24117 oktoberkriget 1
24118 okunnig 3
24119 okunniga 2
24120 okunnighet 6
24121 okunnigt 1
24122 okunskap 1
24123 okuvlig 1
24124 okänd 3
24125 okända 5
24126 okänslig 1
24127 okänsliga 1
24128 okänt 1
24129 olaglig 1
24130 olagliga 3
24131 olagligheter 2
24132 olagligt 5
24133 olet 1
24134 olidliga 1
24135 oligarki 1
24136 oligarkier 1
24137 olik 1
24138 olika 442
24139 olikartade 2
24140 olikhet 1
24141 olikheter 8
24142 olikheterna 4
24143 oliktänkande 1
24144 oliver 3
24145 olivlund 1
24146 olja 11
24147 oljan 7
24148 oljat 1
24149 oljebefraktaren 1
24150 oljeblanka 2
24151 oljebolag 2
24152 oljebolagen 4
24153 oljebolagens 2
24154 oljebolaget 2
24155 oljebälte 7
24156 oljebälten 2
24157 oljebältena 1
24158 oljebältet 7
24159 oljebältets 1
24160 oljeeldningen 1
24161 oljefartyg 4
24162 oljefartygen 1
24163 oljefläckar 1
24164 oljeföroreningar 2
24165 oljeföroreningarna 2
24166 oljeföroreningens 1
24167 oljeindränkta 3
24168 oljeindustrin 1
24169 oljeinkomsterna 1
24170 oljekoka 1
24171 oljekoncernerna 1
24172 oljekontrakt 1
24173 oljelast 1
24174 oljepriser 1
24175 oljeproducenterna 1
24176 oljerester 1
24177 oljeskadefonderna 1
24178 oljeslam 2
24179 oljespill 1
24180 oljestället 1
24181 oljetankbåtar 1
24182 oljetankern 3
24183 oljetankerns 2
24184 oljetankfartyg 2
24185 oljetankfartyget 1
24186 oljetankrar 2
24187 oljetankrarna 1
24188 oljetankrarnas 1
24189 oljetransporter 1
24190 oljetrusterna 1
24191 oljeutsläpp 5
24192 oljeutsläppen 1
24193 oljeutsläppet 1
24194 oljeutvinningsplattformar 1
24195 oljevägen 1
24196 oljig 1
24197 oljiga 2
24198 ologiska 1
24199 olycka 19
24200 olyckan 7
24201 olycklig 5
24202 olyckliga 9
24203 olyckligt 5
24204 olyckligtvis 1
24205 olyckor 20
24206 olyckorna 1
24207 olycksbringande 1
24208 olycksbådande 2
24209 olycksdiger 1
24210 olycksdrabbade 5
24211 olycksfall 1
24212 olycksfallsförsäkringar 1
24213 olycksfåglar 1
24214 olyckshändelse 1
24215 olyckshändelsen 1
24216 olycksrisker 1
24217 olycksriskerna 1
24218 olycksöde 1
24219 olydig 1
24220 olympiska 1
24221 olägenhetslagstiftningarna 1
24222 olämplig 2
24223 olämpliga 3
24224 olämpligt 5
24225 olösligt 1
24226 olösta 3
24227 om 5910
24228 om-ansikte 1
24229 omarbetning 2
24230 ombads 3
24231 ombeds 2
24232 ombesörja 4
24233 ombesörjer 1
24234 ombetts 2
24235 ombonat 1
24236 ombord 10
24237 ombud 2
24238 ombuden 1
24239 ombudsmannen 7
24240 ombudsmannens 8
24241 ombyggnad 1
24242 ombytligt 1
24243 omcentrera 1
24244 omdebatterade 1
24245 omdefiniera 2
24246 omdefinieras 1
24247 omdefiniering 1
24248 omdirigerade 1
24249 omdirigerades 1
24250 omdirigerar 1
24251 omdirigeras 1
24252 omdirigering 1
24253 omdiskuterade 1
24254 omdöme 3
24255 omdömesförmåga 2
24256 omdömesgilla 1
24257 omedelbar 7
24258 omedelbara 5
24259 omedelbart 44
24260 omedgörlig 2
24261 omedveten 2
24262 omedvetet 3
24263 omedvetna 1
24264 omen 1
24265 omfatta 43
24266 omfattade 1
24267 omfattades 3
24268 omfattande 89
24269 omfattar 55
24270 omfattas 33
24271 omfattning 20
24272 omfattningen 8
24273 omflyttning 2
24274 omflyttningar 2
24275 omflyttningen 1
24276 omforma 1
24277 omformulerad 1
24278 omformulerar 1
24279 omformuleras 1
24280 omformulering 2
24281 omfånget 2
24282 omfångsrikt 1
24283 omfördelande 1
24284 omfördelning 5
24285 omfördelningen 2
24286 omförhandlingen 1
24287 omge 1
24288 omger 3
24289 omges 2
24290 omgestaltandet 1
24291 omgift 1
24292 omgivande 3
24293 omgiven 1
24294 omgivet 1
24295 omgivna 1
24296 omgivning 3
24297 omgivningar 2
24298 omgivningarna 1
24299 omgivningen 2
24300 omgruppera 1
24301 omgrupperingar 1
24302 omgående 2
24303 omgång 2
24304 omgångarna 1
24305 omgången 5
24306 omhulda 1
24307 omhändertagandet 1
24308 omintetgör 2
24309 omintetgöra 1
24310 omintetgörs 1
24311 omistlig 1
24312 omklädningsrum 1
24313 omkommit 1
24314 omkostnader 1
24315 omkostnadstäckning 4
24316 omkostnadstäckningen 1
24317 omkramad 1
24318 omkring 91
24319 omkringliggande 1
24320 omkull 1
24321 omkullkastar 1
24322 omlastning 1
24323 omlokaliseringar 3
24324 omlopp 9
24325 omloppsbana 1
24326 ommöblering 1
24327 omnämnande 1
24328 omnämnandena 1
24329 omnämnandet 1
24330 omnämnda 1
24331 omnämnde 1
24332 omnämns 2
24333 omoderna 1
24334 omodernt 2
24335 omogna 1
24336 omoralisk 1
24337 omoraliska 1
24338 omoraliskt 1
24339 omorganisation 1
24340 omorganisationen 7
24341 omorganisera 3
24342 omorganiserar 1
24343 omorganiseras 1
24344 omorganisering 1
24345 omorganiseringen 1
24346 omorientera 1
24347 omotiverat 2
24348 omplacera 1
24349 omplantering 1
24350 omprioritering 1
24351 ompröva 4
24352 omprövar 1
24353 omprövas 2
24354 omprövning 4
24355 omringades 1
24356 område 263
24357 områden 270
24358 områdena 56
24359 områdes 1
24360 områdesbegränsning 1
24361 områdesplaneringen 1
24362 området 222
24363 områdets 1
24364 omröstning 40
24365 omröstningar 9
24366 omröstningarna 5
24367 omröstningen 66
24368 omröstningen.1 1
24369 omröstningsförfarandet 1
24370 omröstningslistan 1
24371 omröstningsregistreringen 1
24372 omröstningsresultaten 1
24373 omsatts 1
24374 omsider 2
24375 omskolning 3
24376 omskrivningar 1
24377 omskärelsen 1
24378 omslag 2
24379 omslaget 1
24380 omsorg 16
24381 omsorgsfulla 1
24382 omsorgsfullt 5
24383 omstridd 3
24384 omstridda 1
24385 omstritt 2
24386 omstrukturera 4
24387 omstrukturering 20
24388 omstruktureringar 7
24389 omstruktureringarna 3
24390 omstruktureringen 2
24391 omstrukturerings- 1
24392 omstruktureringsplan 2
24393 omstruktureringsplaner 1
24394 omstruktureringsåtgärderna 1
24395 omstuvning 1
24396 omställningar 1
24397 omställningen 1
24398 omställningsfasen 1
24399 omständighet 5
24400 omständigheten 3
24401 omständigheter 62
24402 omständigheterna 8
24403 omständliga 2
24404 omsvep 3
24405 omsvängning 2
24406 omsätta 8
24407 omsättas 4
24408 omsätter 1
24409 omsättning 3
24410 omsätts 4
24411 omtalade 4
24412 omtanke 1
24413 omtumlande 1
24414 omtvistad 1
24415 omtvistade 1
24416 omtvistat 1
24417 omvandla 7
24418 omvandlades 1
24419 omvandlar 1
24420 omvandlas 4
24421 omvandlats 2
24422 omvandling 4
24423 omvandlingen 1
24424 omvandlingsprocess 1
24425 omvandlingsprocesser 1
24426 omväg 2
24427 omvägen 1
24428 omvälvande 1
24429 omvälvning 1
24430 omvälvningar 2
24431 omvänd 4
24432 omvända 4
24433 omvänt 7
24434 omvärdera 4
24435 omvärderas 2
24436 omvärdering 2
24437 omvärderingsperioden 1
24438 omvärld 1
24439 omvärlden 2
24440 omväxlande 2
24441 omvårdnad 1
24442 omänsklig 2
24443 omärkliga 1
24444 omärkligt 1
24445 omätliga 1
24446 omålad 1
24447 omöjlig 5
24448 omöjliga 6
24449 omöjligen 2
24450 omöjliggjorde 1
24451 omöjliggör 1
24452 omöjliggörs 2
24453 omöjlighet 1
24454 omöjligheten 1
24455 omöjligt 27
24456 on 2
24457 ond 2
24458 onda 7
24459 ondo 2
24460 ondska 1
24461 ondskan 2
24462 ondskefulla 2
24463 ondskefullt 1
24464 one-stop-shop 1
24465 onekligen 4
24466 online-avtal 1
24467 online-ekonomin 1
24468 onsdag 7
24469 onsdagen 5
24470 onsdags 1
24471 ont 7
24472 onyanserat 1
24473 onödan 1
24474 onödig 6
24475 onödiga 7
24476 onödigt 9
24477 oomkullrunkeliga 1
24478 oomtvistad 1
24479 oordnad 1
24480 oordning 1
24481 oordningen 2
24482 opaler 1
24483 opartisk 1
24484 opartiska 1
24485 opartiskhet 1
24486 opartiskt 4
24487 operahus 1
24488 operan 1
24489 operation 2
24490 operationer 4
24491 operativ 2
24492 operativa 9
24493 operativt 4
24494 operators 1
24495 operatör 1
24496 operatörer 1
24497 operatörerna 2
24498 operera 1
24499 opersonliga 1
24500 opinion 6
24501 opinionen 13
24502 opinioner 2
24503 opinionsbildare 1
24504 opinionsundersökningar 1
24505 oportunidades 1
24506 opp 5
24507 oppe 2
24508 opponera 3
24509 opportunism 1
24510 opportunister 1
24511 opposition 5
24512 oppositionell 1
24513 oppositionen 4
24514 oppositionens 2
24515 oppositionsledaren 1
24516 oppositionspolitikern 1
24517 oppositionstidningar 1
24518 opraktiskt 2
24519 oproportionerliga 2
24520 oproportionerligt 2
24521 optimal 4
24522 optimala 2
24523 optimalt 4
24524 optimera 1
24525 optimeras 1
24526 optimeringen 1
24527 optimism 5
24528 optimistisk 5
24529 optimistiska 2
24530 optimistiskt 4
24531 optioner 3
24532 optionskontrakt 1
24533 optiskt 1
24534 opålitlig 1
24535 orakel 1
24536 orange 2
24537 ord 174
24538 orda 4
24539 ordalag 13
24540 ordalydelsen 2
24541 ordats 1
24542 orden 25
24543 ordentlig 13
24544 ordentliga 1
24545 ordentligt 27
24546 order 6
24547 orders 1
24548 ordet 59
24549 ordförande 203
24550 ordförandebänken 1
24551 ordförandekolleger 1
24552 ordförandeland 1
24553 ordförandelandet 3
24554 ordföranden 25
24555 ordförandena 6
24556 ordförandens 3
24557 ordförandes 1
24558 ordförandeskap 44
24559 ordförandeskapen 2
24560 ordförandeskapens 1
24561 ordförandeskapet 120
24562 ordförandeskapets 31
24563 ordförandeskaps 3
24564 ordförandeskapsprogram 1
24565 ordförandestaten 1
24566 ordinarie 1
24567 ordinär 1
24568 ordlista 1
24569 ordna 6
24570 ordnade 3
24571 ordnandet 1
24572 ordnar 2
24573 ordnas 1
24574 ordnat 2
24575 ordnats 1
24576 ordning 31
24577 ordningar 1
24578 ordningen 13
24579 ordningsfråga 11
24580 ordningsfrågor 2
24581 ordningsfrågorna 2
24582 ordningsföljden 1
24583 ordningsmakt 1
24584 ordre 1
24585 ordrikt 2
24586 ordspråk 1
24587 ordspråket 2
24588 ordvalet 2
24589 ordvrängare 1
24590 ordvändning 1
24591 ordväxlingen 1
24592 orealistisk 2
24593 orealistiska 4
24594 orealistiskt 6
24595 oreda 2
24596 oredan 1
24597 oredlighet 1
24598 oreflekterat 1
24599 oregelbundet 1
24600 oregerliga 1
24601 oreglerade 1
24602 oreglerat 1
24603 oremarkerade 1
24604 organ 49
24605 organen 12
24606 organens 2
24607 organet 3
24608 organisation 25
24609 organisationen 14
24610 organisationens 1
24611 organisationer 63
24612 organisationerna 20
24613 organisationernas 4
24614 organisationers 2
24615 organisations 1
24616 organisationsgraden 1
24617 organisationskapacitet 1
24618 organisationsschema 1
24619 organisationsstruktur 1
24620 organisatoriska 3
24621 organisatoriskt 1
24622 organisera 19
24623 organiserad 4
24624 organiserade 11
24625 organiserades 2
24626 organiserar 6
24627 organiseras 7
24628 organiserats 1
24629 organisering 1
24630 organiskt 1
24631 organism 1
24632 organismer 24
24633 organs 1
24634 orientaler 1
24635 orientaliska 2
24636 orienten 1
24637 orienterad 2
24638 orienterar 1
24639 orienteras 1
24640 orientering 2
24641 orienteringen 1
24642 orienteringsprogrammen 1
24643 originalitet 2
24644 originalspråket 1
24645 originalversionen 3
24646 originella 4
24647 originellt 2
24648 oriktiga 6
24649 oriktigheter 1
24650 oriktigt 2
24651 orimlig 2
24652 orimliga 6
24653 orimligt 3
24654 orkade 2
24655 orkan 1
24656 orkanen 1
24657 orkaner 1
24658 orkester 1
24659 orkestrarnas 1
24660 orm 4
24661 ormen 1
24662 ormens 2
24663 oro 100
24664 oroa 6
24665 oroad 6
24666 oroade 11
24667 oroande 24
24668 oroar 20
24669 oroas 1
24670 orolig 10
24671 oroliga 13
24672 orolige 1
24673 oroligheter 1
24674 oroligt 2
24675 oron 17
24676 orosmoln 2
24677 orosmoment 5
24678 oroväckande 6
24679 orsak 11
24680 orsak-verkanrelationen 1
24681 orsaka 9
24682 orsakade 7
24683 orsakar 10
24684 orsakas 6
24685 orsakat 9
24686 orsakats 7
24687 orsaken 14
24688 orsaker 13
24689 orsakerna 12
24690 orsakssamband 1
24691 orsakssambandet 1
24692 ort 4
24693 orten 4
24694 orter 2
24695 orthomixomicrovirus 1
24696 ortodoxa 2
24697 orubblig 2
24698 orubbliga 2
24699 orwellskt 1
24700 oräkneliga 2
24701 oräkneligt 1
24702 orätt 4
24703 orättfärdiga 1
24704 orättfärdigt 1
24705 orättvis 5
24706 orättvisa 4
24707 orättvisor 7
24708 orättvisorna 3
24709 orättvist 5
24710 orörda 1
24711 orörlig 3
24712 orörlighet 1
24713 orörligt 1
24714 osagt 1
24715 osammanhängande 4
24716 osanna 2
24717 osannolika 3
24718 osar 1
24719 osjälvisk 1
24720 osjälvständiga 1
24721 oskadliga 2
24722 oskakad 1
24723 oskarpa 1
24724 oskiljaktig 1
24725 oskiljaktiga 1
24726 oskriven 1
24727 oskuld 1
24728 oskuldsfull 1
24729 oskuldsfullt 1
24730 oskyldig 2
24731 oskyldiga 2
24732 oskyldigt 1
24733 oslipad 1
24734 osmidig 1
24735 osmältbar 1
24736 osolidariskt 1
24737 oss 1025
24738 ost 2
24739 ostraffade 1
24740 ostron 1
24741 ostronanläggningarna 1
24742 ostronodlare 3
24743 ostronodlarna 2
24744 ostronodling 1
24745 ostronodlingarna 1
24746 ostronodlingarnas 1
24747 ostronodlingen 1
24748 ostrukturerade 1
24749 ostört 1
24750 osv 3
24751 osv. 25
24752 osynlig 2
24753 osynliga 1
24754 osynligt 2
24755 osystematiskt 1
24756 osäker 2
24757 osäkerhet 18
24758 osäkerheten 3
24759 osäkert 2
24760 osäkra 5
24761 osäkrad 1
24762 osäkrare 1
24763 osårbart 1
24764 otacksamma 1
24765 otaliga 4
24766 otillfredsställande 3
24767 otillgängliga 1
24768 otillräcklig 10
24769 otillräckliga 12
24770 otillräcklighet 3
24771 otillräckligheten 1
24772 otillräckligt 10
24773 otillständigt 1
24774 otillåtliga 1
24775 otillåtligt 3
24776 otillåtna 1
24777 otjänlig 1
24778 otjänst 2
24779 otrevligt 1
24780 otrolig 1
24781 otroliga 2
24782 otroligt 3
24783 otrygga 2
24784 otrygghet 2
24785 otryggt 1
24786 otvetydiga 5
24787 otvetydigt 2
24788 otvivelaktig 1
24789 otvivelaktigt 11
24790 otydlig 6
24791 otydliga 3
24792 otydlighet 1
24793 otydligt 4
24794 otyglad 2
24795 otympligt 1
24796 otäckheter 1
24797 otäckt 1
24798 otänkbart 5
24799 otålig 2
24800 otåliga 1
24801 otålighet 2
24802 otåligt 1
24803 ou 2
24804 oumbärlig 2
24805 oumbärliga 2
24806 oumbärligt 4
24807 oundgänglig 1
24808 oundgängliga 4
24809 oundgängligt 1
24810 oundviklig 1
24811 oundvikliga 9
24812 oundvikligen 5
24813 oundvikligt 5
24814 oupphörlig 1
24815 oupphörliga 2
24816 oupplösligt 2
24817 ouppmärksam 1
24818 outbildade 1
24819 outgrundlig 1
24820 outgrundligt 1
24821 outhärdlig 1
24822 outhärdliga 2
24823 outhärdligt 2
24824 outnyttjad 1
24825 outnyttjade 2
24826 outsinlig 1
24827 outsourcing 1
24828 outtalad 1
24829 outtömlig 1
24830 outtömliga 1
24831 outtömligt 1
24832 ovala 1
24833 ovan 5
24834 ovana 1
24835 ovanför 8
24836 ovanifrån 2
24837 ovanlig 2
24838 ovanliga 3
24839 ovanligt 9
24840 ovannämnda 5
24841 ovanpå 6
24842 ovanstående 3
24843 ovederhäftigt 1
24844 over 2
24845 overall 2
24846 overhead-kostnader 1
24847 overkliga 1
24848 overkligt 1
24849 overksam 1
24850 overksamma 1
24851 ovetande 2
24852 oviktiga 1
24853 oviktigt 1
24854 ovilja 3
24855 ovillig 1
24856 ovillkorligen 2
24857 ovisshet 1
24858 oväder 2
24859 ovädren 1
24860 ovädret 1
24861 oväld 1
24862 ovälkomna 1
24863 oväntad 1
24864 oväntade 5
24865 oväntat 6
24866 ovärderlig 2
24867 ovärdig 1
24868 ovärdiga 3
24869 ovärdigt 1
24870 oväsen 1
24871 oväsentligt 1
24872 oändlig 3
24873 oändliga 2
24874 oändlighet 3
24875 oändligheten 1
24876 oändligt 3
24877 oåterkallelig 1
24878 oönskad 2
24879 oönskade 4
24880 oöverlagt 1
24881 oöverskådligt 1
24882 oöverstiglig 3
24883 oöverstigligt 1
24884 oövervinneligt 1
24885 p.17 1
24886 p.g.a. 4
24887 packa 3
24888 packad 1
24889 packat 3
24890 padanska 1
24891 paddlades 1
24892 paket 7
24893 paketet 3
24894 paketsektorn 1
24895 pakten 1
24896 palatsgrindarna 1
24897 palestinier 3
24898 palestinierna 8
24899 palestinsk 2
24900 palestinska 23
24901 palestinskt 2
24902 pall 1
24903 pallen 1
24904 pampig 1
24905 pandemiska 1
24906 paneler 2
24907 panelerna 1
24908 panga 2
24909 panik 3
24910 panikspridning 1
24911 panna 2
24912 pannan 5
24913 pannkaksmakeup 1
24914 pannor 1
24915 panorama 2
24916 panorera 1
24917 pansarattacker 1
24918 pansarvagnar 1
24919 pantomimiskt 1
24920 papegoja 1
24921 papp 3
24922 pappa 7
24923 pappas 2
24924 papper 9
24925 papperet 3
24926 pappersarbete 4
24927 pappersarbetet 2
24928 pappersdokument 1
24929 pappersflagga 1
24930 papperskorgen 1
24931 pappersluntor 1
24932 pappersplaner 1
24933 papperstigrar 1
24934 pappersvaror 1
24935 par 51
24936 paraderade 1
24937 paradigm 3
24938 paradigmskifte 1
24939 paradis 1
24940 paradox 3
24941 paradoxal 3
24942 paradoxala 2
24943 paradoxalt 2
24944 parafraserar 1
24945 paragrafen 1
24946 paragrafrytteriet 1
24947 parallella 9
24948 parallellt 9
24949 paralyseras 1
24950 parameter 1
24951 parametern 1
24952 parametrar 1
24953 parametrarna 1
24954 paramilitära 1
24955 paramilitärt 1
24956 paraply 1
24957 paras 1
24958 parasiter 1
24959 parasoll 1
24960 parcours 1
24961 parece 2
24962 parentes 1
24963 paret 2
24964 parfym 2
24965 paria 1
24966 paritet 1
24967 parité 1
24968 park 2
24969 parken 2
24970 parkens 1
24971 parker 2
24972 parkerad 1
24973 parkerade 2
24974 parkerar 1
24975 parkeringskort 2
24976 parkeringsplatser 1
24977 parlament 135
24978 parlamentariker 14
24979 parlamentarikerna 3
24980 parlamentarisk 11
24981 parlamentariska 19
24982 parlamentariskt 4
24983 parlamentarismen 1
24984 parlamenten 24
24985 parlamentens 2
24986 parlamentet 529
24987 parlamentet- 1
24988 parlamentets 127
24989 parlaments 5
24990 parlamentsbesluten 1
24991 parlamentsbyggnaden 1
24992 parlamentsdebatt 3
24993 parlamentsforum 1
24994 parlamentsgrupp 1
24995 parlamentskolleger 2
24996 parlamentskollegerna 1
24997 parlamentsledamot 16
24998 parlamentsledamoten 3
24999 parlamentsledamöter 29
25000 parlamentsledamöterna 9
25001 parlamentsledamöternas 1
25002 parlamentsnivå 1
25003 parlamentspresidiets 1
25004 parlamentsutskott 3
25005 parlamentsutskotten 1
25006 parlamentsutskottet 1
25007 parmaskinkstunga 1
25008 parningsplatser 1
25009 parodi 1
25010 part 9
25011 parten 3
25012 parter 50
25013 parterna 16
25014 parternas 11
25015 parters 4
25016 parti 52
25017 partiapparaterna 1
25018 partiell 1
25019 partiella 3
25020 partier 24
25021 partierna 13
25022 partiernas 5
25023 partiers 2
25024 partiet 18
25025 partiets 29
25026 partigrupp 3
25027 partigruppen 1
25028 partiintressen 1
25029 partikrati 1
25030 partiledare 1
25031 partimedlems 1
25032 partipolitisk 1
25033 partipolitiska 2
25034 partiprogram 3
25035 partiprogrammet 1
25036 partis 3
25037 partisekreterare 1
25038 partisk 1
25039 partiska 2
25040 partiskt 1
25041 partisplittringens 1
25042 partivänner 1
25043 partner 31
25044 partnern 1
25045 partnerparti 1
25046 partnerrelationen 1
25047 partners 4
25048 partnership 1
25049 partnerskap 41
25050 partnerskapen 3
25051 partnerskapens 1
25052 partnerskapet 8
25053 partnerskapets 2
25054 partnerskaps- 1
25055 partnerskapsavtal 4
25056 partnerskapsavtalen 1
25057 partnerskapsavtalet 4
25058 partnerskapsbidrag 1
25059 partnerskapsformer 1
25060 partnerskapskonceptet 1
25061 partnerskapsländerna 1
25062 partnerskapsmålet 1
25063 partnerskapspolitiken 1
25064 partnerskapsprincipen 3
25065 partnerskapsrådet 1
25066 partnerskapsuppgörelserna 1
25067 partnerstater 1
25068 parts 1
25069 party 1
25070 partyt 1
25071 pas 2
25072 pass 10
25073 passa 10
25074 passade 3
25075 passadvind 1
25076 passage 3
25077 passagerarbuss 1
25078 passagerare 5
25079 passagerarna 7
25080 passagerarnas 1
25081 passagerartransporter 1
25082 passande 10
25083 passar 12
25084 passera 7
25085 passerade 4
25086 passerar 1
25087 passerat 3
25088 passet 1
25089 passion 4
25090 passionerade 1
25091 passionerat 1
25092 passiv 1
25093 passivitet 2
25094 passiviteten 1
25095 passivt 2
25096 passusen 1
25097 pastellmjuka 1
25098 patent 5
25099 patentfrågorna 1
25100 patentmediciner 1
25101 patenträtt 1
25102 patenträttigheterna 1
25103 patentslag 1
25104 paternalistiska 2
25105 paternalistiskt 1
25106 patetisk 1
25107 patetiska 1
25108 patetiskt 1
25109 patient 1
25110 patienter 3
25111 patogen 1
25112 patologiska 1
25113 patriarkalisk 1
25114 patriot 1
25115 patrioters 1
25116 patriotism 1
25117 patrullbåt 1
25118 paus 4
25119 pausen 1
25120 pauser 1
25121 paying 1
25122 peanuts-belopp 1
25123 pedagogiska 2
25124 pedagogiskt 1
25125 pedofilskandaler 1
25126 peka 18
25127 pekade 10
25128 pekar 16
25129 pekat 9
25130 pekfinger 1
25131 pekfingerjingling 1
25132 pelare 10
25133 pelaren 8
25134 pelarna 7
25135 pengar 95
25136 pengarna 33
25137 penna 1
25138 pennan 2
25139 penndrag 1
25140 pennhållare 1
25141 penning- 1
25142 penningdyrkan 1
25143 penningflöden 1
25144 penningflödena 1
25145 penningfurstars 1
25146 penninggirig 1
25147 penningmarknad 1
25148 penningmarknadsinstrument 1
25149 penningmedel 1
25150 penningpolitik 3
25151 penningpolitiken 2
25152 penningpolitisk 1
25153 penningpolitiska 3
25154 penningreferenser 1
25155 penningresurser 1
25156 penningstabilitet 1
25157 penningsummor 1
25158 penningtvätt 4
25159 penningväsendets 1
25160 penny 1
25161 pension 9
25162 pensioner 10
25163 pensioneras 1
25164 pensionerna 8
25165 pensionsbomben 1
25166 pensionsfonder 5
25167 pensionsfondernas 1
25168 pensionsförmånerna 1
25169 pensionsförsäkringarna 1
25170 pensionsmedlen 1
25171 pensionspolitik 1
25172 pensionsrättigheter 1
25173 pensionssystem 2
25174 pensionssystemen 3
25175 pensionssystemens 1
25176 pensionssystemet 2
25177 pensionstidbomb 1
25178 pensionär 3
25179 pensionärer 3
25180 pensionärerna 1
25181 pensionärernas 1
25182 pensionärers 1
25183 per 61
25184 perfekt 12
25185 perfekta 3
25186 pergamentrulle 1
25187 perifera 10
25188 periferin 2
25189 perifert 1
25190 period 32
25191 perioden 60
25192 perioder 5
25193 perioderna 2
25194 periodisk 1
25195 periodiska 15
25196 periodvis 1
25197 perito 1
25198 permanent 7
25199 permanenta 6
25200 perrongen 1
25201 person 36
25202 persona 3
25203 personal 29
25204 personalbrist 1
25205 personaldelen 1
25206 personalen 4
25207 personalens 1
25208 personalförstärkning 1
25209 personalnedskärningar 2
25210 personalnedskärningarna 1
25211 personalpolitik 3
25212 personalpolitiken 1
25213 personalresurser 2
25214 personalresurserna 2
25215 personalsidan 1
25216 personalstrukturen 1
25217 personalutbildning 2
25218 personbil 1
25219 personbyte 1
25220 personell 1
25221 personella 2
25222 personen 2
25223 personer 128
25224 personerna 7
25225 personernas 1
25226 personers 6
25227 personifieras 1
25228 personlandminor 3
25229 personlig 6
25230 personliga 24
25231 personligen 33
25232 personlighet 1
25233 personligheten 1
25234 personligt 4
25235 personne 1
25236 persons 2
25237 persontransporter 1
25238 perspektiv 45
25239 perspektivet 7
25240 peruaner 1
25241 perversas 1
25242 pessimistisk 1
25243 pessimistiskt 1
25244 pest 1
25245 pesten 3
25246 pestens 1
25247 petar 1
25248 petishly 1
25249 petition 1
25250 petroleum 1
25251 pharmaceutiques 1
25252 phtalater 1
25253 piano 1
25254 pickade 1
25255 pickar 1
25256 pickelsburk 1
25257 pickles 1
25258 picknickväska 1
25259 piddlande 1
25260 pigg 1
25261 pikade 1
25262 pikannin 1
25263 pil 1
25264 pilen 2
25265 pilgrimer 2
25266 pilgrimerna 1
25267 piloten 1
25268 piloter 1
25269 pilotfunktion 1
25270 pilotmervärde 1
25271 pilotprogram 2
25272 pilotprojekt 15
25273 pilotstudier 1
25274 pilpilen 1
25275 pincene 1
25276 pinglade 1
25277 pinsam 2
25278 pinsamt 2
25279 pionbusken 1
25280 pionjärer 1
25281 pionjärerna 1
25282 pip 1
25283 pipa 2
25284 pipande 1
25285 pipor 1
25286 pipskägg 1
25287 pir 1
25288 pirat 1
25289 pirater 2
25290 piraternas 1
25291 piratkopiering 1
25292 piratkopior 1
25293 piratversion 1
25294 pirerna 1
25295 piska 1
25296 pivotabellvy 2
25297 pivotdiagramkomponenten 1
25298 pivotdiagramvy 2
25299 pivotdiagramvyns 1
25300 pivottabell 2
25301 pivottabell- 1
25302 pivottabellen 2
25303 pivottabellens 1
25304 pivottabeller 2
25305 pivottabellista 7
25306 pivottabellistan 1
25307 pivottabellistans 1
25308 pivottabellistor 2
25309 pivottabellkomponenten 2
25310 pivottabellvy 5
25311 pivottabellvyer 3
25312 pivottabellvyn 5
25313 pivottabellvyns 1
25314 pivottabelläge 2
25315 pivottabelläget 2
25316 pjäser 1
25317 placera 12
25318 placerad 4
25319 placerade 4
25320 placerades 3
25321 placerar 8
25322 placeras 8
25323 placerat 5
25324 placerats 1
25325 placering 3
25326 placeringen 1
25327 placeringsformerna 1
25328 placeringsmarknaden 2
25329 placeringsmöjligheterna 1
25330 plack 1
25331 pladask 1
25332 pladder 1
25333 plagg 1
25334 plan 41
25335 planekonomiska 1
25336 planen 9
25337 planens 1
25338 planer 32
25339 planera 8
25340 planerad 5
25341 planerade 24
25342 planerades 3
25343 planerande 1
25344 planerar 24
25345 planeras 13
25346 planerat 8
25347 planerats 4
25348 planering 24
25349 planeringen 12
25350 planeringsfasen 2
25351 planeringsskedet 2
25352 planeringsstadiet 1
25353 planerna 7
25354 planet 35
25355 planeten 3
25356 planetens 2
25357 planeter 3
25358 planets 2
25359 plankor 1
25360 plankton 1
25361 planlagda 1
25362 planläggning 1
25363 planlösa 2
25364 planlösningen 1
25365 planlöst 2
25366 plantera 1
25367 plantor 1
25368 plantskolan 1
25369 plast 6
25370 plastbagar 1
25371 plastdisk 1
25372 plasten 1
25373 plastväv 1
25374 plats 91
25375 platsen 17
25376 platser 35
25377 platserna 3
25378 platt 2
25379 platta 4
25380 plattades 1
25381 plattan 2
25382 plattare 1
25383 plattform 1
25384 plattformar 1
25385 plattformsoberoende 1
25386 plattheter 1
25387 plattorna 1
25388 playing 1
25389 plenardebatten 1
25390 plenarkammaren 2
25391 plenarsalen 1
25392 plenarsammanträde 4
25393 plenarsammanträden 1
25394 plenarsammanträdena 1
25395 plenarsammanträdet 7
25396 plenisalen 2
25397 plenum 9
25398 plenumet 2
25399 plikt 11
25400 plikten 2
25401 pliktskyldig 1
25402 plimsollmärket 1
25403 plocka 5
25404 plockade 3
25405 plockats 1
25406 pluggar 1
25407 plumpa 1
25408 plundra 2
25409 plundrare 1
25410 plundras 1
25411 plundring 1
25412 plundringarna 1
25413 plundringen 1
25414 pluralism 1
25415 pluralistiska 4
25416 pluralistiskt 1
25417 plus 5
25418 pluskonto 1
25419 plädera 2
25420 pläderar 5
25421 pläderingen 1
25422 plätt 1
25423 plåga 1
25424 plågade 2
25425 plågar 1
25426 plågas 1
25427 plånboken 2
25428 plånböcker 1
25429 plåt 2
25430 plåtdunk 1
25431 plåtskjul 1
25432 plötslig 3
25433 plötsliga 2
25434 plötsligt 40
25435 poche 1
25436 poena 1
25437 poet 4
25438 poetromantiska 1
25439 poinsettia 1
25440 pojkar 6
25441 pojkarna 1
25442 pojke 12
25443 pojken 9
25444 pojkes 2
25445 poker 1
25446 polacken 1
25447 polacker 1
25448 polackerna 1
25449 polariserat 1
25450 poldermodellen 1
25451 pole 1
25452 polemik 2
25453 polemisk 1
25454 polemiskt 1
25455 polera 1
25456 policy 7
25457 policybeslut 1
25458 policydel 1
25459 policyförslag 1
25460 policyn 2
25461 policyutveckling 1
25462 polis 7
25463 polis- 1
25464 polisakademi 1
25465 polisbevakning 3
25466 polisbyrån 1
25467 polischefen 1
25468 polisen 13
25469 polisenheter 1
25470 polisens 1
25471 poliser 16
25472 polisexperter 1
25473 polisfrågan 1
25474 polisiär 2
25475 polisiära 7
25476 poliskommissarien 1
25477 poliskåren 1
25478 polismyndigheterna 2
25479 polissamarbetet 1
25480 polisstyre 1
25481 polisstyrka 2
25482 polisstyrkan 2
25483 polisstyrkor 1
25484 polisstyrkorna 1
25485 polistjänstemän 2
25486 polisväsendet 1
25487 political 1
25488 politik 317
25489 politiken 111
25490 politikens 7
25491 politiker 27
25492 politikerjargong 1
25493 politikerna 1
25494 politikernas 1
25495 politikers 1
25496 politikområde 4
25497 politikområden 51
25498 politikområdena 6
25499 politikområdenas 2
25500 politiks 2
25501 politiseras 1
25502 politiserat 1
25503 politisk 121
25504 politisk-ekonomiska 1
25505 politiska 376
25506 politiskt 87
25507 pollen 1
25508 polsk 3
25509 polska 3
25510 polske 1
25511 polyaromatisk 1
25512 polycentrisk 1
25513 pompös 1
25514 pompöst 1
25515 pool 1
25516 popularisera 1
25517 populism 1
25518 populismen 1
25519 populistisk 1
25520 populistiska 2
25521 populära 3
25522 porslin 1
25523 porslinsbutik 1
25524 port 1
25525 port-state 2
25526 portarna 1
25527 porten 4
25528 portfölj 4
25529 portföljen 1
25530 portföljer 3
25531 portföljförvaltning 1
25532 portioner 1
25533 portmonnäer 1
25534 portmonnän 1
25535 portokostnad 1
25536 porttelefonen 1
25537 portugis 1
25538 portugisisk 3
25539 portugisiska 126
25540 portugisiske 5
25541 portugisiskt 3
25542 portvin 2
25543 pose 1
25544 posidonia 1
25545 position 12
25546 positionen 3
25547 positioner 6
25548 positiv 68
25549 positiva 72
25550 positivlista 3
25551 positivlistan 1
25552 positivt 81
25553 post 9
25554 posta 1
25555 postala 1
25556 postanställdas 2
25557 postavgifterna 1
25558 postbefordran 1
25559 postbrevbärarna 1
25560 postdirektivet 2
25561 postdistribuerad 1
25562 posten 24
25563 postens 2
25564 poster 11
25565 posterna 4
25566 postföretag 1
25567 postföretagen 4
25568 postförsändelsernas 1
25569 postgången 1
25570 posthandeln 1
25571 posthanteringen 1
25572 postindustriell 1
25573 postindustriella 1
25574 postkoloniala 1
25575 postkontor 13
25576 postkontoren 7
25577 postkontorens 1
25578 postkontoret 2
25579 postkontorsnätverket 1
25580 postkontorstjänster 1
25581 postlåda 1
25582 postmannen 1
25583 postmarknaden 4
25584 postmilitär 1
25585 postmonopolet 1
25586 postområdet 1
25587 postoperatörer 1
25588 postoperatörerna 2
25589 postpolitiken 1
25590 postsektorn 6
25591 postsektorns 2
25592 postservice 2
25593 postsystem 1
25594 posttjänst 2
25595 posttjänstdirektivet 3
25596 posttjänsten 3
25597 posttjänstens 1
25598 posttjänster 29
25599 posttjänsterna 30
25600 posttjänstesektorn 1
25601 posttrafiken 1
25602 postturer 1
25603 posttömningen 1
25604 postutbärare 1
25605 postutbärning 1
25606 postutdelning 2
25607 postutställd 1
25608 postverk 2
25609 postverken 4
25610 postverket 3
25611 postverkets 1
25612 postverksamheten 1
25613 postväsendet 4
25614 potatis 2
25615 potential 13
25616 potentialen 1
25617 potentialer 1
25618 potentiell 3
25619 potentiella 12
25620 potentiellt 3
25621 pottaska 1
25622 poäng 3
25623 poängen 1
25624 poängsystem 4
25625 poängtera 11
25626 poängterar 4
25627 poängterat 3
25628 poängterats 1
25629 ppm 1
25630 prackats 1
25631 practice 1
25632 practice-metoder 1
25633 practices 2
25634 pragmatisk 2
25635 pragmatiska 2
25636 pragmatiskt 2
25637 pragmatism 1
25638 praktexempel 1
25639 praktfull 1
25640 praktfulla 1
25641 praktfullt 1
25642 praktik 3
25643 praktikanter 2
25644 praktiken 35
25645 praktiserar 1
25646 praktiseras 1
25647 praktisk 10
25648 praktiska 33
25649 praktiskt 23
25650 prat 3
25651 prata 20
25652 pratade 4
25653 pratar 5
25654 pratat 2
25655 pratet 1
25656 pratstund 1
25657 praxis 14
25658 praxisen 1
25659 precedensfall 1
25660 precis 99
25661 precisa 5
25662 precisera 5
25663 preciserad 1
25664 preciserade 2
25665 preciserar 3
25666 preciseras 2
25667 preciserat 1
25668 precisering 3
25669 preciseringar 5
25670 precision 6
25671 precist 1
25672 predika 1
25673 predikande 1
25674 prefekt 1
25675 prefektemblem 1
25676 prefekts 1
25677 preferens 2
25678 preferensbehandla 1
25679 preferenser 3
25680 preferensoptionen 1
25681 preferenssystemet 2
25682 prejudicerande 1
25683 prejudikat 6
25684 prelater 1
25685 prelaterna 1
25686 preliminära 5
25687 preliminärt 1
25688 premiss 1
25689 premisser 1
25690 premisserna 1
25691 premiärminister 22
25692 premiärministern 9
25693 premiärministrar 1
25694 premiärministrarna 1
25695 prerogativ 4
25696 prerogativet 1
25697 present 4
25698 presentabla 1
25699 presentation 5
25700 presentationen 5
25701 presentations- 1
25702 presentationsfilen 1
25703 presentationsfiler 1
25704 presentationsformat 3
25705 presentationsinformation 1
25706 presentationsinformationen 1
25707 presenter 3
25708 presentera 22
25709 presenterade 8
25710 presenterades 5
25711 presenterandet 1
25712 presenterar 7
25713 presenteras 13
25714 presenterat 7
25715 presenterats 2
25716 president 29
25717 presidenten 9
25718 presidentens 1
25719 presidenter 1
25720 presidentestraden 1
25721 presidentvalet 1
25722 presidiet 4
25723 presidiets 1
25724 presidium 1
25725 press 8
25726 pressa 3
25727 pressade 5
25728 pressande 1
25729 pressar 2
25730 pressen 15
25731 pressens 2
25732 pressfotografer 1
25733 pressfrihet 5
25734 pressfriheten 2
25735 presskonferens 1
25736 presskonferenser 2
25737 pressmeddelande 1
25738 pressmiddag 1
25739 pressorgan 1
25740 presstjänst 1
25741 prestanda 3
25742 prestation 5
25743 prestationer 2
25744 prestationerna 1
25745 prestationsförmågan 2
25746 prestera 2
25747 presterat 1
25748 preventiv 1
25749 preventiva 1
25750 preventivt 1
25751 prick 1
25752 pricka 1
25753 prickar 2
25754 prickfritt 1
25755 prima 1
25756 primitiva 2
25757 primära 2
25758 primärsektorernas 1
25759 primärt 2
25760 princip 73
25761 principen 98
25762 principer 78
25763 principerna 33
25764 principernas 1
25765 principfast 1
25766 principfrågor 2
25767 principförklaring 1
25768 principförklaringar 1
25769 principiell 1
25770 principiella 3
25771 principiellt 14
25772 principskäl 1
25773 principöverenskommelse 1
25774 prins 1
25775 prinsessan 1
25776 priori 4
25777 prioritera 21
25778 prioriterad 5
25779 prioriterade 16
25780 prioriterades 1
25781 prioriterar 9
25782 prioriteras 16
25783 prioriterat 5
25784 prioritering 8
25785 prioriteringar 31
25786 prioriteringarna 9
25787 prioriteringen 7
25788 prioriteringslistan 1
25789 prioriteringsområden 1
25790 prioriteringsskala 1
25791 prioritet 12
25792 prioriteter 7
25793 prioriteterna 4
25794 priorssäte 1
25795 pris 26
25796 pris- 2
25797 prisa 1
25798 prisade 1
25799 prisas 1
25800 prisats 1
25801 prisberäkningar 1
25802 priser 16
25803 priserna 13
25804 priset 25
25805 prisfastställandet 1
25806 prisgränser 1
25807 prisgränserna 2
25808 prishöjningar 1
25809 prisnivåerna 1
25810 prispolitik 1
25811 prispolitiken 3
25812 prisskillnader 1
25813 prisstabilitet 4
25814 prisstegring 1
25815 prissänkning 1
25816 prissänkningar 1
25817 prissättning 1
25818 prissättningen 2
25819 prisutvecklingen 1
25820 prisökning 2
25821 prisökningen 1
25822 privat 8
25823 privata 56
25824 privatdetektiven 1
25825 privatekonomin 1
25826 privatiseras 1
25827 privatisering 9
25828 privatiseringar 2
25829 privatiseringarna 1
25830 privatiseringen 3
25831 privatiseringens 1
25832 privatlivet 1
25833 privatperson 1
25834 privatpersonen 1
25835 privatpersoner 2
25836 privatsfär 1
25837 privilege 2
25838 privilegier 3
25839 privilegiera 1
25840 privilegierade 2
25841 privilegiet 1
25842 privilegium 5
25843 priviligierade 1
25844 proaktiv 3
25845 problem 369
25846 problematik 1
25847 problematiken 5
25848 problematisk 2
25849 problematiska 1
25850 problematiskt 2
25851 problemen 70
25852 problemens 2
25853 problemet 120
25854 problemets 3
25855 problemlista 1
25856 problemområden 1
25857 problemområdena 3
25858 procedur 3
25859 proceduren 1
25860 procedurer 3
25861 procedurreglerna 1
25862 procent 277
25863 procentandel 2
25864 procentandelarna 1
25865 procenten 3
25866 procents 3
25867 procentsats 3
25868 procentsatsen 1
25869 procentsatser 2
25870 procentsiffror 1
25871 procenttal 3
25872 procenttalet 1
25873 procenttecken 1
25874 procentuellt 1
25875 process 62
25876 processen 48
25877 processens 1
25878 processer 15
25879 processerna 4
25880 processfrågor 2
25881 procession 1
25882 processregler 1
25883 processrättens 1
25884 processuell 1
25885 processuella 4
25886 procès 1
25887 producent 3
25888 producentansvar 3
25889 producentansvaret 3
25890 producenten 6
25891 producentens 2
25892 producenter 11
25893 producenterna 6
25894 producentländerna 1
25895 producera 10
25896 producerade 4
25897 producerar 4
25898 produceras 4
25899 producerat 3
25900 producerats 1
25901 produkt 18
25902 produkten 7
25903 produktens 1
25904 produkter 43
25905 produkterna 4
25906 produkternas 4
25907 produktinnovationer 1
25908 produktion 14
25909 produktionen 5
25910 produktioner 2
25911 produktionsanläggningar 1
25912 produktionsform 1
25913 produktionsföretag 1
25914 produktionskedjan 1
25915 produktionskostnad 1
25916 produktionskostnaderna 2
25917 produktionsled 1
25918 produktionsmedlen 1
25919 produktionsmetod 1
25920 produktionsmetoder 1
25921 produktionsmodell 1
25922 produktionsnedgången 1
25923 produktionsprocessen 1
25924 produktionsresurser 1
25925 produktionssektor 1
25926 produktionssystem 1
25927 produktionsverksamhet 1
25928 produktiv 4
25929 produktiva 8
25930 produktivitet 6
25931 produktiviteten 6
25932 produktivitetsmarginaler 1
25933 produktivitetsstegring 1
25934 produktivitetsvinster 2
25935 produktivitetsvinsterna 1
25936 produktivt 3
25937 produkts 3
25938 professionalism 2
25939 professionell 1
25940 professionella 4
25941 professor 12
25942 profeten 1
25943 profil 3
25944 profilen 1
25945 profilera 1
25946 profilerad 1
25947 profilerat 1
25948 profiterar 1
25949 profylaktisk 1
25950 prognos 2
25951 prognoserna 1
25952 program 232
25953 programansvariga 1
25954 programdokument 1
25955 programförklaring 2
25956 programinitiativen 1
25957 programinriktning 1
25958 programmatiskt 2
25959 programmen 53
25960 programmerar 1
25961 programmeringsspråk 1
25962 programmet 90
25963 programmets 5
25964 programmässiga 2
25965 programmål 1
25966 programperioden 4
25967 programplanering 4
25968 programplaneringen 3
25969 programplaneringsdokument 1
25970 programplaneringsperiod 1
25971 programplaneringsperioden 7
25972 programpunkt 1
25973 programrundan 1
25974 programs 1
25975 programutformningen 1
25976 programvaror 2
25977 programverksamhet 1
25978 progressiv 4
25979 progressiva 1
25980 progressivt 2
25981 prohibition 2
25982 projekt 150
25983 projektadministration 2
25984 projekten 26
25985 projektens 4
25986 projektet 26
25987 projektets 1
25988 projektförslagen 1
25989 projektil 1
25990 projektion 1
25991 projektledningen 2
25992 projektresultat 1
25993 projekts 3
25994 projektvalet 1
25995 proklamera 2
25996 promenad 2
25997 promenaden 1
25998 promenader 2
25999 promenera 2
26000 promenerade 3
26001 promille 1
26002 prompt 1
26003 pronazistiskt 1
26004 propaganda 9
26005 propagandakampanj 1
26006 propagandaskyltar 1
26007 propagera 1
26008 propagerat 2
26009 proportion 6
26010 proportionalitet 1
26011 proportionalitetsprincipen 1
26012 proportionalitetsprinciperna 1
26013 proportionella 1
26014 proportionellt 2
26015 proportioner 2
26016 proportionerliga 1
26017 proppar 1
26018 propuesta 2
26019 prosaiska 1
26020 prospekt 3
26021 prostituerade 2
26022 prostitution 2
26023 prostitutionen 1
26024 proteininnehåll 1
26025 proteinkornspåse 1
26026 protektionism 6
26027 protektionistisk 1
26028 protektionistiska 2
26029 protest 6
26030 protestaktioner 1
26031 protestanter 1
26032 protestantiska 2
26033 protestantiskt 1
26034 protesten 1
26035 protester 7
26036 protestera 2
26037 protesterade 3
26038 protesterar 5
26039 protesterat 2
26040 protestljuden 1
26041 protokoll 14
26042 protokollen 7
26043 protokollet 33
26044 prov 22
26045 prova 1
26046 provanställda 1
26047 provet 1
26048 provins 3
26049 provinsen 4
26050 provinser 1
26051 provinserna 1
26052 provisorisk 2
26053 provisoriska 4
26054 provkandidaterna 1
26055 provkarta 1
26056 provocerande 1
26057 provokation 1
26058 provokationer 1
26059 provunderlag 1
26060 prydd 1
26061 prydligt 1
26062 prydnad 1
26063 prydnadssak 1
26064 prygla 1
26065 pryglades 1
26066 prägel 4
26067 prägeln 2
26068 prägla 3
26069 präglad 5
26070 präglade 3
26071 präglades 1
26072 präglar 2
26073 präglas 7
26074 präglat 1
26075 präglats 3
26076 pråmarna 1
26077 préparez 1
26078 pröva 4
26079 prövade 2
26080 prövar 1
26081 prövas 3
26082 prövats 1
26083 prövning 6
26084 prövningar 3
26085 prövningarna 1
26086 prövoår 1
26087 psalmer 1
26088 pseudo- 1
26089 psykiska 1
26090 psykiskt 1
26091 psykologiska 2
26092 psykologiskt 1
26093 pubar 2
26094 public 1
26095 publicera 1
26096 publicerade 1
26097 publicerades 2
26098 publiceras 1
26099 publicering 1
26100 publicitet 1
26101 publik 2
26102 publiken 1
26103 pudding 2
26104 puertoricansk 1
26105 puffade 1
26106 puls 2
26107 pulserar 1
26108 pulvret 1
26109 pumpa 1
26110 pumpas 4
26111 pund 7
26112 punga 1
26113 pungslagna 1
26114 punkt 227
26115 punkten 84
26116 punkter 100
26117 punkterna 16
26118 punktlig 1
26119 punktligt 1
26120 punkts 1
26121 punktskattepliktiga 1
26122 punktskatter 11
26123 punktskattesats 1
26124 punktskattesatser 1
26125 punktskattesatserna 1
26126 pures 1
26127 puritanska 1
26128 purpurröda 1
26129 pussel 2
26130 pusselbit 1
26131 pusslet 1
26132 putande 1
26133 putsade 2
26134 putsmedel 1
26135 putstrasa 1
26136 pyjamas 1
26137 pyjamasbyxor 1
26138 pyjamasen 2
26139 pyramidisk 1
26140 pälsar 1
26141 pälsverk 1
26142 pärla 1
26143 pärlband 1
26144 pärlbroderier 1
26145 pärlor 2
26146 pärmen 1
26147 päron 1
26148 på 6478
26149 påbjuder 1
26150 påbjudet 1
26151 påbörja 4
26152 påbörjade 3
26153 påbörjades 3
26154 påbörjar 1
26155 påbörjas 3
26156 påbörjat 8
26157 påbörjats 3
26158 pådrag 1
26159 pådrivandet 1
26160 pådyvlas 1
26161 påfallande 3
26162 påfrestande 1
26163 påfrestning 2
26164 påfrestningar 1
26165 påfrestningarnas 1
26166 påfyllning 1
26167 påföljande 2
26168 påföljd 2
26169 påföljden 1
26170 påföljder 3
26171 påföljderna 2
26172 påförde 1
26173 pågick 8
26174 pågå 4
26175 pågående 23
26176 pågår 33
26177 pågått 3
26178 påkalla 1
26179 påkallar 1
26180 påkommen 1
26181 påkopplad 1
26182 pålagor 3
26183 pålar 1
26184 pålitlig 3
26185 pålitliga 2
26186 pålitlighet 1
26187 pålitligt 1
26188 pålägga 1
26189 påläggas 1
26190 påminda 1
26191 påminde 7
26192 påminna 85
26193 påminnande 1
26194 påminnas 2
26195 påminnelse 2
26196 påminner 28
26197 påmint 3
26198 påpeka 59
26199 påpekade 22
26200 påpekades 2
26201 påpekande 8
26202 påpekanden 9
26203 påpekandet 1
26204 påpekar 17
26205 påpekas 5
26206 påpekat 29
26207 påpekats 8
26208 påsen 1
26209 påsk 1
26210 påskynda 7
26211 påskyndade 1
26212 påskyndande 1
26213 påskyndar 1
26214 påskyndas 4
26215 påstod 1
26216 påstods 1
26217 påstridiga 1
26218 påstå 17
26219 påstådd 1
26220 påstående 6
26221 påståenden 3
26222 påståendena 1
26223 påståendet 3
26224 påstår 13
26225 påstås 6
26226 påståtts 2
26227 påstötning 1
26228 påta 1
26229 påtaglig 4
26230 påtagliga 7
26231 påtagligen 1
26232 påtagligt 6
26233 påtala 3
26234 påtalade 2
26235 påtalar 1
26236 påtalat 3
26237 påtalats 5
26238 påtryckning 1
26239 påtryckningar 19
26240 påtryckningarna 2
26241 påtryckningsgrupper 2
26242 påtryckningskampanj 1
26243 påtryckningsmedel 4
26244 påtryckningssanktioner 1
26245 påträffades 1
26246 påträffas 1
26247 påtvinga 3
26248 påtvingad 2
26249 påtvingade 3
26250 påtvingar 1
26251 påtvingas 2
26252 påtvingats 1
26253 påven 2
26254 påverka 27
26255 påverkade 1
26256 påverkan 13
26257 påverkar 40
26258 påverkas 17
26259 påverkat 6
26260 påverkats 8
26261 påvisades 1
26262 påvisar 2
26263 påvisas 1
26264 påvisat 4
26265 påvisats 1
26266 påvisbart 1
26267 pöbelhop 1
26268 qua 3
26269 quality 1
26270 que 1
26271 quidditch 1
26272 quidditchlag 1
26273 quo 3
26274 quota-hoping 1
26275 quoth 1
26276 r 1
26277 rabatt 2
26278 rabatterna 1
26279 rabbi 1
26280 rabbin 1
26281 racerkvast 1
26282 rad 74
26283 rad- 4
26284 raden 4
26285 rader 5
26286 radera 1
26287 raderna 3
26288 radfält 2
26289 radikal 7
26290 radikala 10
26291 radikalernas 1
26292 radikalisering 1
26293 radikalt 9
26294 radio 1
26295 radio- 4
26296 radioaktiva 1
26297 radioaktivt 1
26298 radioamatörfrågan 1
26299 radioklassrum 1
26300 radiologiska 2
26301 radion 4
26302 radioutsändningar 1
26303 radområdet 1
26304 raffinaderier 2
26305 raffinaderiägarna 1
26306 raggiga 1
26307 raiden 2
26308 raisons 1
26309 rak 4
26310 raka 8
26311 rakade 1
26312 rakblad 1
26313 rakbladsskarpa 1
26314 raketanfall 1
26315 raketerna 1
26316 rakryggade 1
26317 raksträcka 1
26318 rakt 14
26319 ram 41
26320 ramar 9
26321 ramarna 6
26322 ramavtal 4
26323 ramavtalet 2
26324 rambeslut 17
26325 rambeslutet 5
26326 rambestämmelser 2
26327 ramdirektiv 10
26328 ramdirektivet 7
26329 ramen 173
26330 ramförslaget 3
26331 ramkonventionen 1
26332 ramlade 4
26333 ramlagstiftning 1
26334 ramlat 1
26335 rammar 1
26336 rampen 1
26337 rampljus 1
26338 rampljuset 1
26339 ramprogram 4
26340 ramprogrammen 1
26341 ramprogrammet 10
26342 ramverk 2
26343 ramvillkor 3
26344 ramvillkoren 2
26345 randområde 1
26346 randområden 9
26347 randområdena 20
26348 randområdet 1
26349 randregioner 1
26350 rang 1
26351 rangordningen 1
26352 rann 3
26353 rannsakande 1
26354 rannsakar 1
26355 rapid 2
26356 rapning 1
26357 rapphöna 1
26358 rappningen 1
26359 rapport 108
26360 rapport.xml 1
26361 rapporten 55
26362 rapportens 4
26363 rapporter 31
26364 rapportera 8
26365 rapporterade 1
26366 rapporterades 1
26367 rapporterar 1
26368 rapporteras 2
26369 rapporterat 2
26370 rapporterats 1
26371 rapportering 5
26372 rapporterna 6
26373 rapportsiffror 1
26374 ras 6
26375 rasade 2
26376 rasande 4
26377 rasat 1
26378 raser 1
26379 rasera 2
26380 raseri 1
26381 rashatet 1
26382 rasisistiska 1
26383 rasism 27
26384 rasismen 5
26385 rasist 1
26386 rasisterna 1
26387 rasistisk 3
26388 rasistiska 18
26389 rasistiskt 5
26390 raskt 2
26391 rasmässig 1
26392 rasslade 2
26393 rast 1
26394 rastillhörighet 1
26395 rastlös 1
26396 rastlösa 2
26397 ratar 1
26398 ratificera 2
26399 ratificerad 1
26400 ratificerade 1
26401 ratificerades 1
26402 ratificerar 4
26403 ratificeras 1
26404 ratificerat 7
26405 ratificerats 2
26406 ratificering 2
26407 ratificeringen 3
26408 ratificeringsförfarandet 1
26409 ratificeringshandlingar 1
26410 ratificeringsprocessen 2
26411 rating 2
26412 rationalisera 5
26413 rationaliserad 1
26414 rationaliserar 1
26415 rationalisering 3
26416 rationaliseringen 1
26417 rationaliseringseffekterna 1
26418 rationell 5
26419 rationella 2
26420 rationellt 5
26421 ratten 1
26422 raucous 1
26423 ravin 1
26424 razzia 2
26425 razzior 1
26426 re-admission 1
26427 reaction 2
26428 reagera 24
26429 reagerade 2
26430 reagerar 7
26431 reagerat 4
26432 reaktion 16
26433 reaktioner 7
26434 reaktionerna 2
26435 reaktionära 1
26436 reaktionärerna 1
26437 reaktionärt 1
26438 reaktorer 8
26439 reaktorhaveri 1
26440 realinkomsten 1
26441 realism 1
26442 realismen 1
26443 realistisk 4
26444 realistiska 8
26445 realistiskt 10
26446 realitet 2
26447 realiteten 11
26448 realiteter 1
26449 realpolitiska 1
26450 realtid 1
26451 rebellerna 2
26452 recept 1
26453 reciprocal 1
26454 recirkulation 1
26455 recognised 1
26456 recovering 1
26457 recycling 1
26458 red 2
26459 reda 28
26460 redaktionella 2
26461 redaktörerna 1
26462 redan 515
26463 redare 1
26464 redares 1
26465 redarna 1
26466 redarnas 1
26467 redas 3
26468 rederi 1
26469 rederier 1
26470 rederiernas 1
26471 rederiet 2
26472 redigera 3
26473 redigerar 3
26474 redlighet 1
26475 redo 9
26476 redogjorde 2
26477 redogjort 4
26478 redogör 2
26479 redogöra 7
26480 redogörelse 5
26481 redogörelsen 1
26482 redogörelser 6
26483 redogörs 1
26484 redovisa 8
26485 redovisade 1
26486 redovisas 1
26487 redovisat 3
26488 redovisats 1
26489 redovisning 3
26490 redovisningskalkylerna 1
26491 redovisningsrubriker 1
26492 redovisningsskyldighet 1
26493 redskap 10
26494 reducera 4
26495 reducerar 1
26496 reduceras 6
26497 reducerat 3
26498 reducerats 1
26499 reducering 2
26500 reduceringen 1
26501 reell 8
26502 reella 8
26503 reellt 2
26504 referensbelopp 3
26505 referensbeloppen 1
26506 referensbibliotek 1
26507 referensen 6
26508 referenser 4
26509 referensfil 1
26510 referensfilen 2
26511 referenspunkt 3
26512 referensram 3
26513 referensramar 2
26514 referensramarna 2
26515 referera 1
26516 refererade 4
26517 refererar 4
26518 refereras 1
26519 reflektera 7
26520 reflektion 2
26521 reflektioner 1
26522 reflektionsarbete 3
26523 reflektionsarbeten 1
26524 reflektionslinje 1
26525 reflektionsplan 1
26526 reflex 1
26527 reflexion 1
26528 reflexionen 1
26529 reflexioner 1
26530 reform 61
26531 reform- 1
26532 reformansträngningar 1
26533 reformarbete 3
26534 reformarbetet 1
26535 reformatorn 1
26536 reformen 29
26537 reformens 6
26538 reformer 48
26539 reformera 14
26540 reformerade 1
26541 reformerar 3
26542 reformeras 6
26543 reformering 12
26544 reformeringen 11
26545 reformeringsmotor 1
26546 reformerna 19
26547 reformförfarande 1
26548 reformförslag 2
26549 reformförslagen 1
26550 reforminstrument 1
26551 reformister 1
26552 reformistisk 1
26553 reformistiska 11
26554 reformpaket 1
26555 reformprocess 4
26556 reformprocessen 7
26557 reformprogram 3
26558 reformprojektet 1
26559 reformsträvanden 1
26560 reformstämpel 1
26561 reformvilja 1
26562 reformvänlig 1
26563 reformvänliga 1
26564 reformåtgärder 1
26565 refuse 1
26566 regel 14
26567 regelbrott 1
26568 regelbunden 4
26569 regelbundenheten 1
26570 regelbundet 21
26571 regelbundna 6
26572 regellös 1
26573 regelmässig 1
26574 regelmässigt 2
26575 regeln 11
26576 regelrätt 1
26577 regelrätta 1
26578 regelsystem 1
26579 regelsystemet 1
26580 regelverk 22
26581 regelverken 1
26582 regelverket 9
26583 regera 1
26584 regerande 4
26585 regerandet 1
26586 regerar 1
26587 regerat 1
26588 regering 87
26589 regeringar 61
26590 regeringarna 41
26591 regeringarnas 7
26592 regeringars 2
26593 regeringen 120
26594 regeringens 20
26595 regerings 3
26596 regeringsbildning 1
26597 regeringsbildningen 9
26598 regeringschef 2
26599 regeringschefer 5
26600 regeringscheferna 9
26601 regeringschefernas 3
26602 regeringsfilosofin 1
26603 regeringsfunktioner 1
26604 regeringsföreträdare 1
26605 regeringsförfarande 1
26606 regeringsförhandlingarna 2
26607 regeringsförklaringen 1
26608 regeringskoalition 2
26609 regeringskoalitionens 1
26610 regeringskonferens 36
26611 regeringskonferensen 122
26612 regeringskonferensens 17
26613 regeringskonferenser 2
26614 regeringskritiker 1
26615 regeringslösningen 1
26616 regeringsmedlemmar 1
26617 regeringsmedlemmarna 1
26618 regeringsmedlemmars 1
26619 regeringsnivå 2
26620 regeringsorgan 1
26621 regeringsorganisationer 1
26622 regeringspartiet 4
26623 regeringsprogram 2
26624 regeringssamarbetets 1
26625 regeringssamarbetsnivå 1
26626 regeringsstrukturen 1
26627 regeringstjänstemän 1
26628 regeringsverksamheten 1
26629 regi 1
26630 regim 7
26631 regimen 9
26632 regimens 2
26633 regimer 4
26634 regimerna 1
26635 region 59
26636 regional 32
26637 regional- 1
26638 regionala 122
26639 regionalisering 1
26640 regionalister 1
26641 regionalplanering 1
26642 regionalplaneringspolitiken 1
26643 regionalpolitik 55
26644 regionalpolitiken 11
26645 regionalpolitikens 2
26646 regionalpolitiska 3
26647 regionalpresident 2
26648 regionalstöd 2
26649 regionalstödet 1
26650 regionalt 13
26651 regionen 73
26652 regionens 6
26653 regioner 145
26654 regionerna 83
26655 regionernas 10
26656 regioners 4
26657 regionnät 1
26658 register 10
26659 registrera 4
26660 registrerad 4
26661 registrerade 2
26662 registrerades 1
26663 registrerar 3
26664 registreras 3
26665 registrerat 1
26666 registrerats 1
26667 registrering 1
26668 registreringen 1
26669 registret 2
26670 regler 111
26671 reglera 16
26672 reglerad 2
26673 reglerade 6
26674 reglerande 3
26675 reglerandet 1
26676 reglerar 10
26677 regleras 14
26678 reglerat 2
26679 reglerats 2
26680 reglering 26
26681 regleringar 3
26682 regleringen 11
26683 regleringsförfarandet 1
26684 regleringskommitté 1
26685 reglerna 43
26686 reglernas 1
26687 regn 4
26688 regna 1
26689 regnade 1
26690 regnar 1
26691 regnbågsringar 1
26692 regndroppsdiamanter 1
26693 regnen 1
26694 regnet 2
26695 regnfloderna 1
26696 regnvatten 1
26697 regressiva 1
26698 reguljära 1
26699 rehabilitering 1
26700 rehabiliteringsprogram 1
26701 rejäl 1
26702 rejäla 3
26703 rejält 6
26704 reklam 6
26705 reklam- 1
26706 reklamdirektör 1
26707 reklamman 1
26708 reklamploj 1
26709 reklamvärldens 1
26710 rekognosceringsturer 1
26711 rekommendation 17
26712 rekommendationen 10
26713 rekommendationer 26
26714 rekommendationerna 19
26715 rekommendera 6
26716 rekommenderade 5
26717 rekommenderades 1
26718 rekommenderar 15
26719 rekommenderas 6
26720 rekommenderat 4
26721 rekonstruktion 2
26722 rekonstruktionsplan 1
26723 rekord 4
26724 rekordlåg 1
26725 rekordsnabb 1
26726 rekordtid 1
26727 rekreationslandskapet 1
26728 rekrytera 1
26729 rekryteringen 1
26730 rekryteringsmetoder 1
26731 rektor 1
26732 relaterade 3
26733 relateras 1
26734 relaterat 1
26735 relation 6
26736 relationen 1
26737 relationer 12
26738 relationerna 9
26739 relativ 6
26740 relativa 2
26741 relativisera 1
26742 relativt 20
26743 relegera 1
26744 relevansen 1
26745 relevant 19
26746 relevanta 17
26747 reliable 1
26748 religion 7
26749 religionsanhängare 1
26750 religiös 2
26751 religiösa 3
26752 religiöst 2
26753 reliken 1
26754 reliker 2
26755 relikerna 1
26756 relikers 1
26757 remiss 1
26758 remora 1
26759 remoran 1
26760 ren 28
26761 rena 24
26762 renar 1
26763 renare 6
26764 renas 1
26765 rengör 1
26766 rengöring 1
26767 rengöringen 1
26768 rengöringskrämer 1
26769 renhet 1
26770 rening 1
26771 reningsstationer 1
26772 reningsverk 2
26773 renligare 1
26774 renovera 1
26775 renoverar 1
26776 renovering 1
26777 renoveringen 1
26778 rensa 6
26779 rensar 1
26780 rensas 1
26781 rensat 2
26782 renskurat 1
26783 rensning 9
26784 rensningen 5
26785 rent 73
26786 rentav 8
26787 rentvättade 1
26788 renässans 1
26789 repade 1
26790 reparationerna 2
26791 reparera 6
26792 reparerat 1
26793 repet 1
26794 repknutar 1
26795 replikerna 1
26796 reportern 1
26797 representant 21
26798 representanten 17
26799 representantens 5
26800 representanter 4
26801 representanthuset 1
26802 representation 10
26803 representationen 2
26804 representationerna 1
26805 representativ 1
26806 representativa 6
26807 representativitet 3
26808 representativt 5
26809 representerad 1
26810 representerade 3
26811 representerar 2
26812 representerat 1
26813 repression 1
26814 repressiva 1
26815 reproduktion 1
26816 reproduktionen 1
26817 reproduktiva 2
26818 reprulle 1
26819 republik 1
26820 republikanerna 4
26821 republikansk 1
26822 republikanska 1
26823 republiken 29
26824 republikens 6
26825 republikerna 2
26826 requis 2
26827 requérant 2
26828 resa 22
26829 resan 1
26830 resande 1
26831 resandet 1
26832 resans 1
26833 researrangörer 1
26834 researrangörernas 2
26835 resejournal 1
26836 resenärer 2
26837 reser 7
26838 reserv 3
26839 reservation 2
26840 reservationer 7
26841 reservationslöst 1
26842 reserven 1
26843 reserver 3
26844 reservera 1
26845 reserverad 1
26846 reserverade 4
26847 reserveras 1
26848 reserverats 1
26849 reservoarpenna 1
26850 reservoarpennor 1
26851 reservtrupper 1
26852 reseslitna 1
26853 residens 1
26854 residuer 1
26855 resignera 1
26856 resklar 1
26857 resning 1
26858 resolut 2
26859 resolution 117
26860 resolutionen 81
26861 resolutionen.)Talmannen 1
26862 resolutionens 2
26863 resolutioner 26
26864 resolutionerna 6
26865 resolutionsförslag 37
26866 resolutionsförslagen 2
26867 resolutionsförslaget 14
26868 resolutionsförslagets 1
26869 resolutionstext 1
26870 resonanslåda 1
26871 resonemang 7
26872 resonemangen 2
26873 resonemanget 1
26874 resonera 1
26875 resonerade 2
26876 resonliga 1
26877 resor 4
26878 resource 1
26879 resp. 2
26880 respekt 79
26881 respektabel 1
26882 respektabelt 1
26883 respektabilitet 2
26884 respekten 34
26885 respektera 30
26886 respekterade 2
26887 respekterar 31
26888 respekteras 28
26889 respekterat 1
26890 respektfull 1
26891 respektingivande 2
26892 respektive 44
26893 respons 4
26894 responsibilise 1
26895 rest 5
26896 rest-Jugoslavien 1
26897 restaurang 2
26898 restaurangen 1
26899 restaurangförbunden 1
26900 restaureringsarbetena 1
26901 reste 10
26902 resten 20
26903 rester 1
26904 resterande 4
26905 resterna 2
26906 restriktion 1
26907 restriktioner 2
26908 restriktionerna 3
26909 restriktiv 1
26910 restriktiva 1
26911 restriktivt 1
26912 rests 1
26913 restvara 1
26914 restämnen 1
26915 resultant 1
26916 resultat 146
26917 resultaten 37
26918 resultatet 43
26919 resultatinriktad 1
26920 resultatlista 1
26921 resultattavla 6
26922 resultattavlan 1
26923 resultatöversikt 4
26924 resultatöversikten 2
26925 resultera 1
26926 resulterade 3
26927 resulterar 8
26928 resulterat 5
26929 resurs 13
26930 resursbristen 1
26931 resursen 3
26932 resurser 115
26933 resurserna 36
26934 resursernas 2
26935 resursfrågor 1
26936 resursförbrukningskostnaderna 1
26937 resursfördelning 2
26938 resursförvaltning 1
26939 resurskrävande 1
26940 resursproblem 1
26941 resursslöseri 1
26942 resurstilldelning 1
26943 resväska 2
26944 resårer 1
26945 reta 1
26946 retar 1
26947 retirera 1
26948 retorik 12
26949 retroaktiv 1
26950 retroaktiva 3
26951 retroaktivitet 3
26952 retroaktiviteten 1
26953 retroaktivt 5
26954 retrospektiv 1
26955 reträtt 4
26956 returnerar 3
26957 rev 1
26958 revben 3
26959 revidera 8
26960 reviderade 3
26961 revideras 4
26962 revidering 17
26963 revideringar 1
26964 revideringen 10
26965 revideringsklausul 1
26966 revideringsklausulen 1
26967 revirstrider 1
26968 revision 6
26969 revisionen 1
26970 revisionsarbetskommittén 1
26971 revisionsarbetskommittés 1
26972 revisionsenheten 1
26973 revisionsfunktioner 1
26974 revisionsförklaring 1
26975 revisionsförklaringen 1
26976 revisionsroller 1
26977 revisionsrätten 13
26978 revisionsrättens 6
26979 revisionssystem 2
26980 revisionstjänst 2
26981 revisionstjänsten 2
26982 revisionsuppföljning 1
26983 revisorns 1
26984 revolution 6
26985 revolutionen 3
26986 revolutioner 1
26987 revolutionslandet 1
26988 revolutionsregeringens 1
26989 revolutionär 4
26990 revolutionära 3
26991 revolver 1
26992 ribban 1
26993 rida 2
26994 ridande 1
26995 riddare 3
26996 rider 2
26997 ridning 1
26998 ridå 1
26999 ridån 1
27000 riggade 1
27001 rights 1
27002 rigiditeten 1
27003 rigorös 1
27004 rigorösa 3
27005 rigoröst 4
27006 rik 5
27007 rika 20
27008 rikare 3
27009 rikaste 5
27010 rikedom 8
27011 rikedomar 8
27012 rikedomarna 3
27013 rikedomen 6
27014 riket 2
27015 riklig 5
27016 rikligt 1
27017 riksdagen 1
27018 riksdagens 1
27019 riksdagsledamöter 1
27020 rikt 4
27021 rikta 27
27022 riktad 4
27023 riktade 15
27024 riktades 1
27025 riktar 12
27026 riktas 10
27027 riktat 3
27028 riktats 2
27029 riktig 24
27030 riktiga 8
27031 riktige 1
27032 riktigt 83
27033 riktlinje 2
27034 riktlinjen 2
27035 riktlinjer 86
27036 riktlinjerna 42
27037 riktlinjernas 3
27038 riktning 61
27039 riktningar 1
27040 riktningarna 2
27041 riktningen 16
27042 riktpunkter 2
27043 rimlig 12
27044 rimliga 14
27045 rimligare 1
27046 rimligen 2
27047 rimligt 16
27048 rimligtvis 1
27049 rimmar 1
27050 ring 2
27051 ringa 12
27052 ringakta 1
27053 ringde 8
27054 ringen 1
27055 ringer 8
27056 ringklockan 1
27057 ringlade 1
27058 ringt 1
27059 rinner 1
27060 ris 2
27061 risk 36
27062 riskabel 3
27063 riskanalys 3
27064 riskavfall 1
27065 riskbedömning 3
27066 riskbedömningen 1
27067 risken 39
27068 risker 32
27069 riskera 7
27070 riskerade 1
27071 riskerar 43
27072 riskerna 17
27073 riskexponering 1
27074 riskfaktor 1
27075 riskfritt 1
27076 riskfylld 2
27077 riskfyllda 4
27078 riskfyllt 2
27079 riskförebyggande 2
27080 riskhantering 5
27081 riskhanteringsfunktion 1
27082 riskkapital 6
27083 riskkommunikation 2
27084 risknivå 1
27085 riskspridning 1
27086 riskspridningsprincipen 1
27087 riskspridningsregler 2
27088 risktagande 2
27089 risktagarna 1
27090 riskuppgifterna 1
27091 riskutvecklingen 1
27092 riskvilligt 1
27093 riskvärdering 3
27094 riskzonen 2
27095 riste 1
27096 ritat 1
27097 ritualbärare 1
27098 ritualen 1
27099 rituell 1
27100 rituella 1
27101 riva 1
27102 rivalen 1
27103 rivs 1
27104 ro 7
27105 roade 5
27106 roar 2
27107 roat 2
27108 robusta 1
27109 rock 2
27110 rocken 1
27111 rockfickan 1
27112 rockskört 1
27113 roder 2
27114 rodnaden 1
27115 rodret 1
27116 roffa 1
27117 rofylld 1
27118 rogivande 1
27119 roliga 1
27120 roligt 12
27121 roll 221
27122 rollen 12
27123 roller 4
27124 roman 1
27125 romaner 1
27126 romantik 1
27127 romantiken 1
27128 romantiska 1
27129 romarna 2
27130 romarnas 1
27131 romer 6
27132 romerbefolkningen 1
27133 romergruppen 1
27134 romerna 2
27135 romernas 1
27136 ropa 2
27137 ropade 7
27138 ropande 1
27139 ropar 4
27140 ropet 2
27141 ros 3
27142 rosa 5
27143 rosafärgad 1
27144 rosenröd 1
27145 rosenrött 1
27146 rosig 1
27147 rosor 1
27148 rosorna 2
27149 rostade 3
27150 rostar 1
27151 rostat 2
27152 rostbildning 1
27153 rostig 2
27154 rostiga 1
27155 rota 1
27156 rotade 2
27157 rotat 1
27158 rotation 1
27159 rotelement 1
27160 rotelementet 1
27161 roten 1
27162 rotsystem 1
27163 rott 1
27164 round 1
27165 rovfiske 1
27166 rubba 1
27167 rubbar 1
27168 rubbas 1
27169 rubbat 1
27170 rubbats 1
27171 rubbningarna 1
27172 rubrik 14
27173 rubriken 3
27174 rubriker 2
27175 rubrikerna 1
27176 ruelse 1
27177 ruffig 1
27178 ruffiga 1
27179 rufsiga 1
27180 rufsigt 1
27181 rugbybrede 1
27182 ruin 2
27183 ruiner 2
27184 ruinerad 1
27185 ruineras 1
27186 ruinerna 1
27187 ruljangsen 1
27188 rullade 3
27189 rullande 1
27190 rullar 4
27191 rullat 2
27192 rullats 1
27193 rullstol 1
27194 rullstolen 1
27195 rullstolsburna 1
27196 rum 142
27197 rumlade 1
27198 rummel 1
27199 rummet 24
27200 rumänsk 1
27201 rumänska 4
27202 rund 1
27203 runda 8
27204 rundabordskonferens 1
27205 rundan 3
27206 rundor 2
27207 rundresa 3
27208 rundresan 1
27209 rundtur 1
27210 runt 62
27211 runtom 2
27212 rusa 3
27213 rusade 11
27214 rusande 1
27215 rusar 4
27216 rusat 1
27217 ruskig 1
27218 rusningen 1
27219 rusningstiden 1
27220 rusta 2
27221 rustad 2
27222 rustningsproblemets 1
27223 rutan 1
27224 rutig 1
27225 rutin 2
27226 rutinen 2
27227 rutiner 12
27228 rutinerna 3
27229 rutinmässiga 2
27230 rutmönster 1
27231 rutnät 1
27232 rutnätets 2
27233 ruttna 3
27234 ruttnade 2
27235 ruttnande 1
27236 ruvade 3
27237 ruvande 2
27238 ryck 1
27239 rycka 2
27240 rycker 2
27241 ryckig 1
27242 ryckigt 1
27243 ryckte 7
27244 rycktes 1
27245 ryckts 1
27246 rygg 6
27247 rygga 2
27248 ryggar 1
27249 ryggen 10
27250 ryggmusklerna 1
27251 ryggrad 3
27252 ryggraden 1
27253 ryktas 1
27254 ryktbarhet 1
27255 rykte 7
27256 rykten 3
27257 ryktena 1
27258 rymde 2
27259 rymden 7
27260 rymdmonster 1
27261 rymdtid 2
27262 rymdåldern 1
27263 rymma 2
27264 rymmer 2
27265 ryms 1
27266 rynkor 1
27267 rysk 2
27268 ryska 17
27269 ryske 9
27270 rysligt 1
27271 rysning 3
27272 ryssar 1
27273 ryssarna 7
27274 ryste 1
27275 rytm 3
27276 rytmiskt 1
27277 ryttarna 1
27278 räcka 16
27279 räcker 59
27280 räckhåll 4
27281 räcks 1
27282 räckte 13
27283 räckvidd 6
27284 rädd 15
27285 rädda 30
27286 räddade 2
27287 räddades 1
27288 räddande 1
27289 räddar 2
27290 räddas 1
27291 räddat 2
27292 räddats 1
27293 räddning 3
27294 räddningen 2
27295 räddningshelikoptrar 2
27296 räddningsnivåer 1
27297 räddningstjänst 1
27298 räddningstjänster 1
27299 rädsla 10
27300 rädslan 5
27301 räkenskap 2
27302 räkenskaper 1
27303 räkenskaperna 7
27304 räkenskapsansvariga 1
27305 räkenskapssystemet 1
27306 räkenskapsår 1
27307 räkna 26
27308 räknade 3
27309 räknar 39
27310 räknas 7
27311 räknat 8
27312 räknats 1
27313 räkneexempel 1
27314 räkning 31
27315 räkningar 1
27316 räkningen 2
27317 räls 1
27318 räntan 1
27319 räntehöjning 1
27320 ränteintäkter 1
27321 ränteutgifter 1
27322 räntor 1
27323 räntorna 1
27324 rät 1
27325 räta 1
27326 rätade 1
27327 rätas 1
27328 rätt 286
27329 rätta 74
27330 rättade 1
27331 rättades 1
27332 rättan 1
27333 rättar 1
27334 rättas 3
27335 rättats 2
27336 rättegång 6
27337 rättegångar 2
27338 rättegången 1
27339 rättegångsprocesser 1
27340 rätteligen 2
27341 rättelse 1
27342 rätten 72
27343 rättens 1
27344 rättfram 2
27345 rättframt 2
27346 rättfärdiga 6
27347 rättfärdigande 1
27348 rättfärdiganden 1
27349 rättfärdigandet 1
27350 rättfärdigar 4
27351 rättfärdigas 2
27352 rättfärdigat 1
27353 rättfärdigt 1
27354 rättighet 23
27355 rättigheten 1
27356 rättigheter 276
27357 rättigheterna 174
27358 rättigheternas 5
27359 rättigheters 1
27360 rättighetsinnehavarna 2
27361 rättighetsstadgor 1
27362 rättmätig 2
27363 rättmätiga 2
27364 rättmätigt 2
27365 rättrogna 1
27366 rättrådigheten 1
27367 rätts- 1
27368 rättsakt 4
27369 rättsakter 3
27370 rättsdefinition 1
27371 rättsförluster 1
27372 rättshjälp 20
27373 rättshjälpen 4
27374 rättsinniga 1
27375 rättsinstanser 2
27376 rättsinstanserna 1
27377 rättskaffens 2
27378 rättskipning 7
27379 rättskipningssystemet 1
27380 rättskultur 1
27381 rättskulturen 1
27382 rättslig 55
27383 rättsliga 164
27384 rättsligt 37
27385 rättsläget 3
27386 rättsområde 2
27387 rättsordning 1
27388 rättsordningen 2
27389 rättsosäkerhet 2
27390 rättspraxis 3
27391 rättsprincip 1
27392 rättsprinciper 1
27393 rättsprocess 1
27394 rättsprocessen 2
27395 rättsregler 1
27396 rättsreglerna 1
27397 rättssamarbetet 1
27398 rättssekreterare 1
27399 rättsskipande 3
27400 rättsskipning 2
27401 rättsskipningen 2
27402 rättsskydd 1
27403 rättsskyddsområdet 1
27404 rättsstat 5
27405 rättsstaten 4
27406 rättsstatens 2
27407 rättsstatliga 1
27408 rättsstatlighet 2
27409 rättsstatsprincip 1
27410 rättsstatsprincipen 2
27411 rättsstatus 1
27412 rättsstödet 1
27413 rättssystem 17
27414 rättssystemen 8
27415 rättssystemet 7
27416 rättssäkerhet 15
27417 rättssäkerheten 8
27418 rättstillämpningen 1
27419 rättstjänst 1
27420 rättstjänsten 1
27421 rättstraditionen 1
27422 rättstraditioner 2
27423 rättsuppfattningen 1
27424 rättsutskottet 1
27425 rättsutskottets 1
27426 rättsväsen 1
27427 rättsväsende 4
27428 rättsväsendet 3
27429 rätttsliga 1
27430 rättvis 28
27431 rättvisa 85
27432 rättvisan 10
27433 rättvisans 2
27434 rättvisare 2
27435 rättvisebehov 1
27436 rättvisefrågor 1
27437 rättvisekriterier 1
27438 rättvist 29
27439 rättänkande 1
27440 rå 1
27441 råa 1
27442 råare 1
27443 råd 40
27444 råda 24
27445 rådande 8
27446 rådde 8
27447 rådens 2
27448 råder 71
27449 rådet 506
27450 rådets 269
27451 rådfråga 3
27452 rådfrågade 1
27453 rådfrågades 2
27454 rådfrågar 2
27455 rådfrågat 2
27456 rådfrågats 2
27457 rådfrågningar 1
27458 rådfrågningsprocessen 1
27459 rådgivande 14
27460 rådgivare 5
27461 rådgivarna 1
27462 rådgivarnas 1
27463 rådgivning 7
27464 rådgivningen 1
27465 rådgivningsnätverk 1
27466 rådgivningsverksamhet 1
27467 rådgör 1
27468 rådighet 1
27469 råds 2
27470 rådsbeslut 1
27471 rådsbeslutet 1
27472 rådsförsamlingar 1
27473 rådsgruppen 1
27474 rådslag 3
27475 rådsledamöterna 1
27476 rådsmedlemmar 1
27477 rådsministrar 1
27478 rådsmötena 1
27479 rådsmötet 9
27480 rådsordförande 55
27481 rådsordföranden 18
27482 rådsordförandens 3
27483 rådsordförandeskapet 3
27484 rådsordförandeskapets 1
27485 rådsrepresentanternas 1
27486 rådsresolution 1
27487 rådstoppmötet 1
27488 rågata 1
27489 råkade 5
27490 råkar 4
27491 råkat 2
27492 råmaterial 3
27493 råmärken 1
27494 rånade 1
27495 rånares 1
27496 rånkupp 1
27497 råolja 3
27498 råskinn 1
27499 rått 4
27500 råtta 2
27501 råttan 1
27502 råttor 1
27503 råvara 1
27504 råvaror 1
27505 råvarorna 1
27506 råvaruproducenter 1
27507 référendaire 1
27508 röd 9
27509 röda 21
27510 rödgröna 1
27511 rödhårig 1
27512 rödklädda 1
27513 rödrutig 1
27514 rödvin 1
27515 rödögda 1
27516 rök 2
27517 röka 2
27518 röken 1
27519 röker 2
27520 rökgrå 1
27521 rökmoln 1
27522 rökningen 1
27523 rökpuffar 1
27524 rökridåer 1
27525 rökte 5
27526 rönt 1
27527 rönte 1
27528 rör 115
27529 röra 19
27530 röran 1
27531 rörande 64
27532 röras 1
27533 rörde 15
27534 rörelse 12
27535 rörelsehindrade 1
27536 rörelsen 3
27537 rörelser 8
27538 rörelserna 1
27539 rören 1
27540 rörig 1
27541 rörigt 3
27542 rörlig 2
27543 rörliga 4
27544 rörlighet 30
27545 rörligheten 18
27546 rört 5
27547 röst 45
27548 rösta 112
27549 röstade 37
27550 röstades 3
27551 röstar 37
27552 röstas 4
27553 röstat 40
27554 röstats 1
27555 rösten 6
27556 röster 20
27557 rösterna 2
27558 röstförklaring 7
27559 röstförklaringar 1
27560 röstförklaringarna 1
27561 röstkapacitet 1
27562 röstlista 1
27563 röstresultat 1
27564 rösträtt 4
27565 rösträtten 3
27566 röstsystem 2
27567 röstsystemet 2
27568 röstsystemsfråga 1
27569 röstviktning 3
27570 röta 1
27571 rött 9
27572 rötter 5
27573 rötterna 2
27574 röv 1
27575 rövats 1
27576 s 3
27577 s'il 1
27578 s. 1
27579 s.16 1
27580 s.k. 16
27581 sa 123
27582 sabbaten 1
27583 sabeltandad 1
27584 sadaterna 1
27585 sade 266
27586 sades 3
27587 safety-protokollet 1
27588 sagan 1
27589 sagda 1
27590 sagt 160
27591 sagts 32
27592 sak 118
27593 sak- 3
27594 sak-om-faktisk 1
27595 saken 38
27596 sakens 4
27597 saker 116
27598 sakerna 7
27599 sakernas 2
27600 sakfrågan 3
27601 sakfrågor 2
27602 sakförhållanden 1
27603 sakförhållandena 1
27604 sakinnehållet 1
27605 sakkunnig 1
27606 sakkunniga 6
27607 sakkunskap 4
27608 sakkunskapen 1
27609 sakkännedom 2
27610 saklig 1
27611 sakliga 2
27612 sakligt 1
27613 sakna 1
27614 saknade 9
27615 saknaden 1
27616 saknades 3
27617 saknar 34
27618 saknas 58
27619 saknat 2
27620 saknats 1
27621 sakområden 1
27622 sakområdet 1
27623 sakproblem 1
27624 sakta 16
27625 sakupplysning 1
27626 sal 1
27627 salen 2
27628 salinarbetare 1
27629 salladsblad 1
27630 salong 2
27631 saltdofter 1
27632 saltvatten 1
27633 salu 2
27634 saluföra 2
27635 saluförande 1
27636 saluförandet 1
27637 saluförde 1
27638 saluföringen 3
27639 saluföringsfrågorna 1
27640 saluföringskostnaderna 1
27641 saluförs 2
27642 salutant 1
27643 samarbeta 27
27644 samarbetar 12
27645 samarbetat 3
27646 samarbete 169
27647 samarbetet 86
27648 samarbetets 3
27649 samarbets- 3
27650 samarbetsanda 4
27651 samarbetsavtal 4
27652 samarbetsavtalet 3
27653 samarbetsbetonat 1
27654 samarbetskapacitet 1
27655 samarbetsklimat 1
27656 samarbetskommittén 1
27657 samarbetsländerna 1
27658 samarbetsmodell 1
27659 samarbetsområden 1
27660 samarbetsområdena 2
27661 samarbetsorganisation 1
27662 samarbetspartner 1
27663 samarbetspolitik 5
27664 samarbetspolitiken 5
27665 samarbetsprincipen 1
27666 samarbetsprocess 1
27667 samarbetsprogram 1
27668 samarbetsprojekt 3
27669 samarbetsprojekten 1
27670 samarbetsramen 1
27671 samarbetsstrategi 1
27672 samarbetssätt 1
27673 samarbetsutveckling 1
27674 samarbetsvilja 1
27675 samarbetsvilliga 1
27676 samband 139
27677 sambanden 2
27678 sambandet 4
27679 samexistens 7
27680 samexistensen 1
27681 samfinansierades 1
27682 samfinansieras 1
27683 samfinansiering 2
27684 samfinansieringen 1
27685 samfund 1
27686 samfunden 2
27687 samfundet 12
27688 samfundets 3
27689 samförstånd 21
27690 samförståndspolitik 1
27691 samhälle 50
27692 samhällelig 2
27693 samhälleliga 3
27694 samhällen 33
27695 samhällena 5
27696 samhälles 4
27697 samhället 79
27698 samhällets 15
27699 samhällsaktörer 1
27700 samhällsansvar 1
27701 samhällsekonomin 1
27702 samhällsekonomisk 1
27703 samhällsekonomiska 3
27704 samhällsfaktor 1
27705 samhällsfientliga 1
27706 samhällsgrupperna 1
27707 samhällsklasser 1
27708 samhällskostnaderna 1
27709 samhällsliv 2
27710 samhällslivet 1
27711 samhällsmedborgare 1
27712 samhällsmodell 1
27713 samhällsmodellen 3
27714 samhällsomfattande 11
27715 samhällsomgivningen 1
27716 samhällsområden 1
27717 samhällspolitiska 1
27718 samhällsservicen 1
27719 samhällsstöd 1
27720 samhällssystem 1
27721 samhällsteori 1
27722 samhällsvärde 1
27723 samhörande 1
27724 samhörigheten 1
27725 samklang 2
27726 samla 22
27727 samlad 2
27728 samlade 14
27729 samlades 3
27730 samlar 3
27731 samlarfordon 1
27732 samlarmani 1
27733 samlas 7
27734 samlat 10
27735 samlats 5
27736 samlevnad 3
27737 samlevnaden 1
27738 samlevnadsformer 1
27739 samling 7
27740 samlingsplatser 1
27741 samma 300
27742 sammalunda 1
27743 samman 57
27744 sammanbindande 1
27745 sammanblanda 1
27746 sammanblandning 2
27747 sammanboende 1
27748 sammanbrott 1
27749 sammanbunden 1
27750 sammandrabbning 1
27751 sammandrag 1
27752 sammanfalla 1
27753 sammanfallande 1
27754 sammanfallanden 1
27755 sammanfaller 5
27756 sammanfatta 8
27757 sammanfattade 1
27758 sammanfattande 1
27759 sammanfattar 4
27760 sammanfattas 3
27761 sammanfattat 2
27762 sammanfattning 10
27763 sammanfattningar 1
27764 sammanfattningen 1
27765 sammanfattningsvis 6
27766 sammanflätade 2
27767 sammanfogas 1
27768 sammanfogat 1
27769 sammanför 1
27770 sammanföra 5
27771 sammanföras 1
27772 sammanförde 1
27773 sammanhang 85
27774 sammanhangen 2
27775 sammanhanget 50
27776 sammanhopningen 2
27777 sammanhängande 10
27778 sammanhänger 1
27779 sammanhållande 2
27780 sammanhållen 2
27781 sammanhållning 63
27782 sammanhållningen 45
27783 sammanhållningsfonden 1
27784 sammanhållningsländerna 2
27785 sammanhållningspolitik 3
27786 sammanhållningspolitiken 2
27787 sammanhållningspolitikens 2
27788 sammanhållningsprocessen 2
27789 sammanhörande 2
27790 sammanjämka 2
27791 sammanjämkar 1
27792 sammankalla 5
27793 sammankallande 2
27794 sammankallandet 4
27795 sammankallas 1
27796 sammankomst 1
27797 sammankomster 2
27798 sammankomsterna 1
27799 sammankoppla 1
27800 sammankopplade 2
27801 sammanlagd 1
27802 sammanlagda 3
27803 sammanlagt 4
27804 sammanlänka 1
27805 sammanlänkade 1
27806 sammansatt 7
27807 sammansatta 1
27808 sammanslaget 1
27809 sammanslagning 3
27810 sammanslagningar 6
27811 sammanslagningen 4
27812 sammanslagningsvåg 1
27813 sammanslutning 2
27814 sammanslutningar 6
27815 sammanslutningarna 2
27816 sammanslutnings 1
27817 sammansmältningens 1
27818 sammanställa 2
27819 sammanställd 1
27820 sammanställde 1
27821 sammanställer 1
27822 sammanställning 6
27823 sammanställningen 4
27824 sammanställs 1
27825 sammanställt 2
27826 sammanställts 1
27827 sammansvärjning 1
27828 sammansättning 6
27829 sammansättningen 6
27830 sammanträda 3
27831 sammanträdde 1
27832 sammanträde 30
27833 sammanträden 4
27834 sammanträdena 4
27835 sammanträder 4
27836 sammanträdesperiod 7
27837 sammanträdesperioden 2
27838 sammanträdesperiodens 1
27839 sammanträdesperioder 1
27840 sammanträdesperioderna 1
27841 sammanträdesrum 1
27842 sammanträdessessionen 1
27843 sammanträdestakten 1
27844 sammanträdet 25
27845 sammanträdets 1
27846 sammanträffande 1
27847 sammanträffanden 1
27848 sammanträtt 1
27849 sammetsdraperade 1
27850 sammetsstol 1
27851 samordna 26
27852 samordnad 11
27853 samordnade 13
27854 samordnande 2
27855 samordnar 2
27856 samordnare 4
27857 samordnarna 1
27858 samordnas 5
27859 samordnat 3
27860 samordnats 1
27861 samordning 60
27862 samordningen 25
27863 samordningsaspekt 1
27864 samordningsförfarandet 1
27865 samordningsförmåga 1
27866 samordningsmekanismer 1
27867 samordningsmetod 1
27868 samordningsproblem 1
27869 samordningsprocess 1
27870 samordningsstruktur 1
27871 samriskföretag 2
27872 samråd 19
27873 samråda 3
27874 samråden 2
27875 samrådet 2
27876 samrådsakt 1
27877 samrådsarbete 1
27878 samrådsdirektiv 1
27879 samrådsdokumentet 1
27880 samrådsforum 1
27881 samrådsförfarande 1
27882 samrådsförfaranden 1
27883 samrådsförfarandet 1
27884 samrådsförslaget 1
27885 samrådskommittéer 1
27886 samrådsprocess 1
27887 samrådsprocessen 1
27888 samrådsrättigheter 1
27889 samsats 1
27890 samspel 1
27891 samspelet 2
27892 samspråk 1
27893 samstämmig 6
27894 samstämmiga 3
27895 samstämmighet 63
27896 samstämmigheten 21
27897 samstämmighetsobservatorium 1
27898 samstämmighetspolitiken 1
27899 samstämmighetsprocessen 1
27900 samstämmighetsövervakning 1
27901 samstämmigt 7
27902 samstämt 1
27903 samsyn 5
27904 samt 230
27905 samtal 35
27906 samtala 2
27907 samtalande 1
27908 samtalar 1
27909 samtalen 13
27910 samtalet 8
27911 samtalspartner 3
27912 samtalsrundan 1
27913 samtalssvårigheter 1
27914 samtalsämne 1
27915 samtida 2
27916 samtidens 1
27917 samtidighet 1
27918 samtidigt 188
27919 samtliga 91
27920 samtycke 17
27921 samtycker 3
27922 samtyckesförfarandet 2
27923 samtyckt 1
27924 samvarotid 1
27925 samverka 6
27926 samverkan 5
27927 samverkande 1
27928 samverkar 2
27929 samvete 1
27930 samveten 3
27931 samvetet 3
27932 samvetsgranna 1
27933 samvetslös 1
27934 samvetsskäl 1
27935 sandaler 2
27936 sanden 1
27937 sandtag 1
27938 sanera 4
27939 sanerats 1
27940 saneringen 8
27941 saneringsarbete 1
27942 sanitär 2
27943 sanitära 3
27944 sanka 1
27945 sanktion 1
27946 sanktionen 1
27947 sanktioner 29
27948 sanktionera 2
27949 sanktionerad 1
27950 sanktionerna 7
27951 sanktionspolitik 1
27952 sanktionssystem 2
27953 sanktionssystemet 1
27954 sann 2
27955 sanna 3
27956 sannerligen 13
27957 sanning 4
27958 sanningen 13
27959 sanningens 1
27960 sannings- 1
27961 sannolika 2
27962 sannolikhet 5
27963 sannolikheten 1
27964 sannolikhetskalkyl 1
27965 sannolikt 16
27966 sansad 1
27967 sansat 2
27968 sant 47
27969 sargande 1
27970 sarkastisk 1
27971 satellit 2
27972 satelliter 1
27973 satellitteve 1
27974 satellitövervakning 2
27975 satsa 24
27976 satsade 1
27977 satsar 6
27978 satsas 3
27979 satsat 3
27980 satsats 1
27981 satsning 8
27982 satsningar 4
27983 satsningen 3
27984 satt 62
27985 satta 3
27986 satte 29
27987 sattes 5
27988 satts 6
27989 scale 1
27990 scen 1
27991 scenarbetare 1
27992 scenarier 3
27993 scenario 2
27994 scenarior 1
27995 scenariot 2
27996 scenen 5
27997 scener 1
27998 schablonmässiga 1
27999 schablonmässigt 1
28000 schackbräde 1
28001 schema 7
28002 scheman 3
28003 schemat 5
28004 schizofren 1
28005 schweiziska 2
28006 scientifiques 1
28007 scones 1
28008 sconesen 1
28009 scoreboard 1
28010 se 533
28011 securities 2
28012 sedan 363
28013 sedda 1
28014 seder 1
28015 sedlar 2
28016 sedlarna 2
28017 sedligt 1
28018 sedvanliga 3
28019 sedvanor 1
28020 seg 2
28021 segdraget 1
28022 segel 1
28023 segelbara 1
28024 segelfartyg 1
28025 segelleden 1
28026 seger 7
28027 segern 3
28028 segla 5
28029 seglade 4
28030 seglar 14
28031 seglat 1
28032 seglen 2
28033 seglingen 1
28034 segment 1
28035 segra 1
28036 segrat 1
28037 seismisk 1
28038 seismiska 1
28039 sekel 12
28040 sekellång 1
28041 sekellöst 1
28042 sekelskifte 1
28043 sekelskiftet 1
28044 sekelslutet 1
28045 sekler 1
28046 seklerna 1
28047 seklers 1
28048 seklet 2
28049 sekretariat 4
28050 sekretariatet 1
28051 sekreterare 3
28052 sekreteraren 1
28053 sekretess 6
28054 sekretessbelagd 1
28055 sekretessbelagda 3
28056 sekretessbelägga 1
28057 sekretessbelägger 1
28058 sekretessen 1
28059 sekretesshänsynen 1
28060 sekretessstadga 1
28061 sekretion 1
28062 sektion 3
28063 sektionerna 1
28064 sektor 39
28065 sektorer 46
28066 sektorerna 11
28067 sektoriell 3
28068 sektoriella 2
28069 sektorinriktad 2
28070 sektorinriktade 1
28071 sektorintressen 1
28072 sektorn 43
28073 sektorns 10
28074 sektorpolitik 1
28075 sektors 1
28076 sektorsanalys 1
28077 sektorsfråga 1
28078 sektorsinriktat 1
28079 sektorsspecifika 1
28080 sektorsövergripande 2
28081 sekulariserade 1
28082 sekund 4
28083 sekunder 6
28084 sekundärprocesser 1
28085 sekundärrätten 1
28086 sekundärtransvestit 1
28087 seldon 1
28088 selektiv 5
28089 selektiva 6
28090 selektivitet 1
28091 selektivt 8
28092 semantisk 1
28093 semester 8
28094 semesterfirare 1
28095 semesterfirarna 1
28096 semestertider 1
28097 semestra 1
28098 semestrar 1
28099 semestrarna 1
28100 seminarier 1
28101 seminarierna 1
28102 seminariet 1
28103 seminarium 3
28104 sen 18
28105 sena 3
28106 senare 110
28107 senareläggas 2
28108 senareläggning 1
28109 senast 20
28110 senaste 173
28111 senat 2
28112 senaten 2
28113 senator 4
28114 senatorer 1
28115 senfärdig 1
28116 sensibilitet 1
28117 sent 30
28118 sentimentalitet 1
28119 separat 6
28120 separata 8
28121 separatism 1
28122 separerade 2
28123 separerat 1
28124 september 27
28125 ser 262
28126 sera 1
28127 serb 1
28128 serber 16
28129 serberna 4
28130 serbisk 1
28131 serbiska 7
28132 serie 8
28133 seriefält 1
28134 serier 1
28135 seriesläppområde 1
28136 seriös 5
28137 seriösa 6
28138 seriösare 1
28139 seriöst 20
28140 servats 1
28141 servera 3
28142 serverad 1
28143 serverades 1
28144 serverar 1
28145 serveringsfat 1
28146 service 30
28147 serviceföretag 1
28148 servicekort 1
28149 servicekvalitet 2
28150 servicen 15
28151 servicenivå 1
28152 servicens 1
28153 servicenätverk 1
28154 ses 32
28155 session 20
28156 sessionen 20
28157 sessioner 3
28158 sessionerna 1
28159 sessionstiden 1
28160 sessionstjänsten 1
28161 sett 140
28162 setts 1
28163 sex 50
28164 sex- 1
28165 sex-trettio 1
28166 sexismen 1
28167 sexmånadersperiod 3
28168 sextio 2
28169 sextiotalet 4
28170 sextiotusenmannastyrkan 1
28171 sextiotvå 1
28172 sexton 4
28173 sextumskanonerna 2
28174 sexturismen 1
28175 sexuell 2
28176 sexuella 3
28177 sexuellt 2
28178 sexvärt 1
28179 sexårsdag 1
28180 sexårsperiod 1
28181 sfär 2
28182 sfärer 1
28183 shall 1
28184 shamprocks 1
28185 sharing 1
28186 sherry 1
28187 shilling 1
28188 shipping 1
28189 shirt-fronter 1
28190 shorts 2
28191 shownummer 1
28192 si 1
28193 sicilianska 1
28194 sicksackade 1
28195 sida 146
28196 sidan 203
28197 sidans 1
28198 siden 1
28199 sidenklänning 1
28200 sidenträ 1
28201 sidfilnamn.bak.htm 1
28202 sidfot 1
28203 sidfotsektion 1
28204 sidhuvud 1
28205 sidhuvudsektion 1
28206 sidoblick 1
28207 sidoeffekter 1
28208 sidor 28
28209 sidorna 11
28210 siffermässiga 1
28211 siffra 7
28212 siffran 1
28213 siffror 19
28214 siffrorna 13
28215 sig 1792
28216 signal 20
28217 signalen 2
28218 signaler 7
28219 signalerar 2
28220 signerade 1
28221 signerar 1
28222 signerat 1
28223 signifikant 1
28224 signifikativt 1
28225 signum 1
28226 sikt 62
28227 sikta 2
28228 siktade 1
28229 siktar 6
28230 sikte 8
28231 siktet 1
28232 sill 1
28233 sillhuvuden 2
28234 silver 4
28235 silver- 1
28236 silverfärgade 1
28237 silverförvanskningen 1
28238 silvergarnityr 1
28239 silverglänsande 1
28240 silverräv 1
28241 silversiklar 1
28242 silverskimrande 1
28243 silvertråden 1
28244 simma 1
28245 simpel 2
28246 simpla 1
28247 simulatorer 2
28248 sin 639
28249 sina 462
28250 sinad 1
28251 sine 5
28252 singel 1
28253 sinnade 1
28254 sinnat 1
28255 sinne 4
28256 sinnelag 3
28257 sinnen 3
28258 sinnena 1
28259 sinnesrörelse 2
28260 sinnesstämning 1
28261 sinnet 1
28262 sinom 2
28263 sinsemellan 9
28264 sir 3
28265 sist 47
28266 sista 109
28267 siste 2
28268 sistnämnda 11
28269 sistnämndas 1
28270 sistone 1
28271 sitt 369
28272 sitta 15
28273 sittande 2
28274 sittbad 1
28275 sitter 33
28276 sittning 2
28277 situation 131
28278 situationen 176
28279 situationens 6
28280 situationer 30
28281 situationerna 1
28282 sjabbig 1
28283 sjabbiga 1
28284 sjabblar 1
28285 sjok 1
28286 sju 27
28287 sjudande 1
28288 sjuhundra 2
28289 sjuk 12
28290 sjuk- 2
28291 sjuka 4
28292 sjukdom 11
28293 sjukdomar 12
28294 sjukdomen 8
28295 sjukdomens 2
28296 sjukdomsbekämpning 1
28297 sjukdomsskydd 1
28298 sjuke 1
28299 sjukes 1
28300 sjukförsäkring 1
28301 sjukhus 9
28302 sjukhusen 1
28303 sjukhuset 7
28304 sjukhusplatserna 1
28305 sjukligt 2
28306 sjukvård 3
28307 sjukvården 1
28308 sjukvårdens 1
28309 sjukvårds- 1
28310 sjukvårdsanläggningar 1
28311 sjukvårdsbudgeten 1
28312 sjukvårdsfrågorna 1
28313 sjukvårdspolitik 1
28314 sjunde 5
28315 sjunga 3
28316 sjungande 2
28317 sjunger 2
28318 sjunka 10
28319 sjunkande 1
28320 sjunken 1
28321 sjunker 3
28322 sjunkit 10
28323 sjunkna 5
28324 sjutton 2
28325 sjuttonde 1
28326 sjuårsperiod 2
28327 själ 7
28328 själar 2
28329 själen 2
28330 själlösa 1
28331 själv 226
28332 själva 244
28333 självaktning 1
28334 självaste 1
28335 självbedrägeri 1
28336 självbedrägerier 1
28337 självbelåtenhet 1
28338 självbelåtne 1
28339 självbestämmande 6
28340 självbiografi 4
28341 självbärande 2
28342 självdeskriptiva 1
28343 självdispergerad 1
28344 självfallet 7
28345 självförnöjelse 1
28346 självförsörjande 2
28347 självförtroende 1
28348 självförtroendet 1
28349 självförvaltande 1
28350 självförvållade 1
28351 självhjälp 3
28352 självklar 7
28353 självklara 4
28354 självklarhet 6
28355 självklart 49
28356 självkostnadspriser 1
28357 självkänsla 1
28358 självlysande 1
28359 självmant 1
28360 självmedlidande 1
28361 självmord 1
28362 självplågeri 1
28363 självreglerande 1
28364 självrespekt 1
28365 självstympning 1
28366 självstyrande 6
28367 självstyre 2
28368 självstyrelse 3
28369 självstyrelsens 1
28370 självstyrelseorganen 1
28371 självstyret 1
28372 självständig 6
28373 självständiga 8
28374 självständighet 5
28375 självständigheten 1
28376 självständighetsbalen 1
28377 självständighetsceremonin 1
28378 självständighetsdagen 1
28379 självständighetsfesten 2
28380 självständighetsfirandet 2
28381 självständighetsparti 1
28382 självständighetsprocess 1
28383 självständighetsrörelsen 2
28384 självständigt 10
28385 självsäkert 3
28386 självt 22
28387 självtillit 1
28388 självtäkt 1
28389 självuttryck 1
28390 självverkande 1
28391 självändamål 4
28392 sjätte 21
28393 sjättedel 1
28394 sjöar 3
28395 sjöarna 1
28396 sjöcertifikat 1
28397 sjöd 1
28398 sjödugligt 1
28399 sjöfarande 1
28400 sjöfarandes 1
28401 sjöfarten 1
28402 sjöfartens 1
28403 sjöfartsinspektionen 1
28404 sjöfartsmyndigheter 1
28405 sjöfartsområdena 1
28406 sjöfartsorganisationen 2
28407 sjöfartssektorn 3
28408 sjöfolk 1
28409 sjögående 1
28410 sjöman 5
28411 sjömannamässigt 1
28412 sjömannen 1
28413 sjömansbalaklava 1
28414 sjömän 3
28415 sjömännen 3
28416 sjön 11
28417 sjöng 5
28418 sjönk 10
28419 sjöovärdiga 1
28420 sjörätt 1
28421 sjöss 7
28422 sjöstjärnor 1
28423 sjösäkerhet 4
28424 sjösäkerheten 3
28425 sjösättas 1
28426 sjötransport 1
28427 sjötransporten 1
28428 sjötransporter 3
28429 sjötransportsektorn 1
28430 sjövägen 1
28431 sjövärdighetscertifikat 1
28432 ska 55
28433 skada 38
28434 skadad 1
28435 skadade 6
28436 skadades 2
28437 skadan 3
28438 skadar 18
28439 skadas 2
28440 skadat 3
28441 skadats 6
28442 skadeersättning 1
28443 skadeersättningsanspråk 1
28444 skadeglädje 1
28445 skadegörelse 1
28446 skademinskning 1
28447 skadestånd 1
28448 skadeståndsfrågorna 1
28449 skadlig 8
28450 skadliga 18
28451 skadligare 1
28452 skadligaste 1
28453 skadligt 6
28454 skador 40
28455 skadorna 14
28456 skadornas 2
28457 skaffa 20
28458 skaffade 1
28459 skaffar 2
28460 skaffat 3
28461 skaka 2
28462 skakade 8
28463 skakande 1
28464 skakar 2
28465 skakat 3
28466 skakningar 1
28467 skal 2
28468 skala 7
28469 skalan 1
28470 skaldjur 1
28471 skaldjuren 1
28472 skaldjursfisket 1
28473 skall 1904
28474 skalle 1
28475 skallen 1
28476 skallig 2
28477 skalligt 1
28478 skam 7
28479 skamfläck 1
28480 skamlig 3
28481 skamliga 1
28482 skamligt 3
28483 skammen 1
28484 skampålen 3
28485 skandal 8
28486 skandalanklagelserna 1
28487 skandalen 1
28488 skandaler 1
28489 skandalerna 4
28490 skandalös 1
28491 skandalösa 2
28492 skandalöst 5
28493 skapa 298
28494 skapad 1
28495 skapade 9
28496 skapades 6
28497 skapande 7
28498 skapandet 38
28499 skapandets 1
28500 skapar 90
28501 skapare 4
28502 skaparens 1
28503 skaparkraften 1
28504 skapas 44
28505 skapat 22
28506 skapats 20
28507 skapelsen 1
28508 skapelsens 1
28509 skapular 1
28510 skar 3
28511 skara 2
28512 skaran 3
28513 skarp 3
28514 skarpa 4
28515 skarpsinniga 2
28516 skarpt 7
28517 skarv 1
28518 skatt 13
28519 skatta 1
28520 skatte- 2
28521 skatteaspekterna 1
28522 skattebasen 1
28523 skattebestämmelser 1
28524 skattebestämmelserna 1
28525 skattebetalare 10
28526 skattebetalaren 1
28527 skattebetalarna 9
28528 skattebetalarnas 3
28529 skattebördan 1
28530 skatteflykt 1
28531 skattefria 1
28532 skattefrågan 2
28533 skattefrågor 4
28534 skatteförvaltningen 1
28535 skatteförändringar 1
28536 skatteharmonisering 3
28537 skatteharmoniseringen 1
28538 skatteincitament 1
28539 skatteindrivares 1
28540 skatteinkomster 1
28541 skatteinspektörer 1
28542 skattekonkurrens 1
28543 skatteliknande 2
28544 skattelättnader 3
28545 skattemässig 1
28546 skattemässiga 6
28547 skattemässigt 1
28548 skatten 1
28549 skatteområdet 5
28550 skatteparadis 2
28551 skattepengar 2
28552 skattepolitik 3
28553 skattepolitiken 4
28554 skatter 14
28555 skattereform 2
28556 skatteregler 1
28557 skatterna 2
28558 skattesamordning 3
28559 skattesamordningen 1
28560 skattesats 1
28561 skattesatser 1
28562 skattesatserna 1
28563 skattestrukturen 1
28564 skattesystem 2
28565 skattesystemet 4
28566 skattetryck 1
28567 skattetrycket 2
28568 skatteuppgifter 1
28569 skatteändringar 1
28570 skatteåtgärder 1
28571 skattkista 1
28572 skattsedeln 2
28573 ske 95
28574 sked 1
28575 skedd 1
28576 skedde 13
28577 skede 18
28578 skeden 1
28579 skedet 2
28580 sken 8
28581 skenat 1
28582 skenet 1
28583 skenhelighet 1
28584 skenheligt 1
28585 skenorna 1
28586 skepnader 1
28587 skepp 4
28588 skeppare 1
28589 skeppas 1
28590 skeppat 1
28591 skeppen 1
28592 skeppsbrott 1
28593 skeppsbrottet 1
28594 skeppsbyggnad 1
28595 skeppslanternor 1
28596 skeppsredare 2
28597 skeppsredarnas 1
28598 skeppsvarv 1
28599 skeppsvarven 1
28600 skepsis 2
28601 skepticismen 1
28602 skeptiker 1
28603 skeptisk 6
28604 skeptiska 1
28605 skeptiskt 1
28606 sker 115
28607 skett 50
28608 skick 14
28609 skicka 21
28610 skickad 2
28611 skickade 11
28612 skickades 5
28613 skickar 9
28614 skickas 5
28615 skickat 3
28616 skickats 2
28617 skicklig 3
28618 skicklighet 1
28619 skickligt 2
28620 skifta 2
28621 skiftade 1
28622 skiftande 1
28623 skiftning 1
28624 skikt 2
28625 skilda 14
28626 skilde 1
28627 skildes 2
28628 skildra 1
28629 skildrar 2
28630 skildrats 2
28631 skildring 1
28632 skilja 5
28633 skiljaktigheter 1
28634 skiljaktigheterna 1
28635 skiljas 2
28636 skiljedomare 1
28637 skiljedomarna 1
28638 skiljedomsprövning 1
28639 skiljeförfarandena 1
28640 skiljelinjer 1
28641 skiljer 33
28642 skiljt 1
28643 skillnad 27
28644 skillnaden 13
28645 skillnader 36
28646 skillnaderna 31
28647 skilsmässa 2
28648 skilsmässan 1
28649 skimrade 2
28650 skinande 1
28651 skiner 1
28652 skingra 2
28653 skingrades 1
28654 skinkomeletter 1
28655 skinkor 1
28656 skinkstek 1
28657 skipa 2
28658 skipas 3
28659 skir 1
28660 skiss 3
28661 skissar 1
28662 skissera 3
28663 skisserade 1
28664 skisseras 1
28665 skisserat 2
28666 skit 1
28667 skiva 1
28668 skivor 1
28669 skivsuccéerna 1
28670 skivtallriken 1
28671 skjorta 3
28672 skjortan 4
28673 skjul 3
28674 skjulet 1
28675 skjuta 18
28676 skjutas 7
28677 skjutberedd 1
28678 skjuter 9
28679 skjutit 1
28680 skjutits 6
28681 skjuts 9
28682 skjutvapen 1
28683 sko 4
28684 skog 5
28685 skogar 20
28686 skogarna 13
28687 skogarnas 3
28688 skogen 6
28689 skogklädda 1
28690 skogrikedomar 1
28691 skogsarbetarna 1
28692 skogsavverkningen 1
28693 skogsbefolkningens 1
28694 skogsberoende 1
28695 skogsbolagens 1
28696 skogsbruk 1
28697 skogsbrukarna 1
28698 skogsbruket 6
28699 skogsfastighet 1
28700 skogsförordningen 1
28701 skogskommuner 1
28702 skogskornell 1
28703 skogslagar 1
28704 skogsodlingsmaterial 1
28705 skogsområden 1
28706 skogsområdena 1
28707 skogspolitik 1
28708 skogssektorn 3
28709 skogssektorns 1
28710 skogsskövlingen 1
28711 skogsutrustning 1
28712 skogsägaren 2
28713 skoja 1
28714 skojigt 1
28715 skola 8
28716 skolan 14
28717 skolans 1
28718 skolböcker 1
28719 skolelev 1
28720 skolelever 1
28721 skolflicka 1
28722 skolflickor 1
28723 skolformelböcker 1
28724 skollista 1
28725 skolläraraktig 1
28726 skolmaten 1
28727 skolor 4
28728 skolorna 1
28729 skolprefekter 1
28730 skolsalar 1
28731 skolundervisning 1
28732 skolåret 1
28733 skon 1
28734 skona 2
28735 skonar 1
28736 skonas 1
28737 skoningslös 1
28738 skoningslöst 1
28739 skor 1
28740 skorna 1
28741 skorpiga 1
28742 skorsten 2
28743 skorstenar 1
28744 skorstenen 1
28745 skotsk 3
28746 skotska 14
28747 skotske 1
28748 skotskt 1
28749 skotten 1
28750 skramlade 1
28751 skrammel 1
28752 skrap 1
28753 skrapa 2
28754 skrapie 11
28755 skrapningar 1
28756 skratt 13
28757 skratta 3
28758 skrattade 15
28759 skrattande 2
28760 skrattas 1
28761 skrattet 1
28762 skrattretande 1
28763 skrattspegel 1
28764 skrek 4
28765 skrev 19
28766 skrevs 4
28767 skriade 1
28768 skriande 1
28769 skribenter 1
28770 skrider 1
28771 skriftlig 5
28772 skriftliga 5
28773 skriftligen 8
28774 skriftligt 8
28775 skrik 4
28776 skrika 2
28777 skrikande 1
28778 skrin 1
28779 skriv 1
28780 skriva 28
28781 skrivas 1
28782 skrivberedd 1
28783 skrivbord 3
28784 skrivbordet 1
28785 skrivbordsliv 1
28786 skrivbordsstolen 1
28787 skrivbordsutvärdering 1
28788 skrivelse 10
28789 skrivelsen 3
28790 skrivelser 2
28791 skriven 2
28792 skriver 9
28793 skrivet 4
28794 skrivfel 1
28795 skrivit 21
28796 skrivits 2
28797 skrivna 4
28798 skrivningar 1
28799 skrivskyddat 1
28800 skrot 1
28801 skrota 1
28802 skrotade 2
28803 skrotar 2
28804 skrotas 5
28805 skrotfärdigt 1
28806 skrotning 5
28807 skrotningen 2
28808 skrotningsföretag 2
28809 skrotningskostnaden 1
28810 skrotningskostnaderna 1
28811 skrotningsprocesserna 1
28812 skrotningssystem 1
28813 skrov 5
28814 skrovet 2
28815 skrovkonstruktionens 1
28816 skrovsidan 1
28817 skrubb 1
28818 skrubben 2
28819 skrumpnad 1
28820 skrumpnade 1
28821 skrupelfria 2
28822 skrupler 1
28823 skrupulös 1
28824 skrynklade 1
28825 skrynkliga 2
28826 skryt 1
28827 skryta 3
28828 skryter 1
28829 skrytsamt 1
28830 skräck 2
28831 skräckens 1
28832 skräckinjagande 1
28833 skräckscenarior 1
28834 skräckslagen 1
28835 skräckväldet 1
28836 skräddarsydda 1
28837 skräddarsytt 1
28838 skräll 1
28839 skrällande 1
28840 skrämd 1
28841 skrämde 2
28842 skrämma 1
28843 skrämmande 3
28844 skrämmas 1
28845 skrämmer 2
28846 skräms 1
28847 skräp 2
28848 skräpet 3
28849 skräpiga 1
28850 skräpuppsamlarsyssla 1
28851 skugga 6
28852 skuggad 4
28853 skuggan 5
28854 skuggboxningen 1
28855 skuggig 2
28856 skuggor 3
28857 skuggorna 3
28858 skuggparlament 1
28859 skuld 2
28860 skuldavskrivning 1
28861 skuldbelägger 1
28862 skuldbörda 1
28863 skuldbördan 1
28864 skulden 4
28865 skulder 4
28866 skulderna 1
28867 skuldfullt 1
28868 skuldkvittning 1
28869 skuldmedvetet 1
28870 skuldmedvetna 1
28871 skuldnivåerna 1
28872 skuldnivån 1
28873 skuldsanering 1
28874 skuldsättning 2
28875 skuldsättningen 1
28876 skuldutvecklingen 1
28877 skull 39
28878 skulle 1652
28879 skumma 1
28880 skummjölksblått 1
28881 skumpade 1
28882 skumrasket 1
28883 skumögda 1
28884 skurarna 1
28885 skurits 1
28886 skurkar 1
28887 skurkarna 1
28888 skuta 1
28889 skutan 2
28890 skutt 1
28891 skutta 1
28892 skuttande 1
28893 skvaller 1
28894 skvalpade 1
28895 skydd 86
28896 skydda 79
28897 skyddad 1
28898 skyddade 6
28899 skyddande 1
28900 skyddar 12
28901 skyddas 11
28902 skyddat 3
28903 skyddet 49
28904 skydds- 1
28905 skyddsbestämmelser 1
28906 skyddsbestämmelserna 2
28907 skyddsgallren 1
28908 skyddsklausuler 1
28909 skyddslingar 1
28910 skyddslösa 1
28911 skyddsnivå 5
28912 skyddsnivån 4
28913 skyddsnät 2
28914 skyddsnäten 1
28915 skyddsområde 6
28916 skyddsområdet 4
28917 skyddsrum 1
28918 skyddsstyrka 1
28919 skyddssystemen 1
28920 skyddstullar 1
28921 skyddstullarna 1
28922 skyddsvärn 1
28923 skyddsåtgärder 1
28924 skyfall 1
28925 skyfallen 1
28926 skyfflade 1
28927 skygga 1
28928 skygghet 1
28929 skyhöga 1
28930 skyhögt 1
28931 skyla 3
28932 skyldig 14
28933 skyldiga 27
28934 skyldighet 26
28935 skyldigheten 6
28936 skyldigheter 21
28937 skyldigt 2
28938 skylla 1
28939 skyllas 1
28940 skyller 1
28941 skylten 2
28942 skyltfönster 2
28943 skyltfönstret 1
28944 skyltning 1
28945 skymda 1
28946 skymma 2
28947 skymningen 3
28948 skymningsljus 1
28949 skymt 2
28950 skymta 1
28951 skymtade 3
28952 skymtande 2
28953 skymtat 2
28954 skymts 1
28955 skymundan 1
28956 skyn 1
28957 skynda 8
28958 skyndade 6
28959 skyndar 3
28960 skyndsamhet 1
28961 skyndsamt 6
28962 skyttevärn 1
28963 skägget 5
28964 skäggprydd 1
28965 skäggstubb 2
28966 skäl 100
28967 skälen 11
28968 skälet 25
28969 skälig 4
28970 skäliga 4
28971 skäligen 1
28972 skäligt 3
28973 skämdes 1
28974 skämma 2
28975 skämmas 4
28976 skäms 2
28977 skämt 2
28978 skämtade 1
28979 skämtar 1
28980 skämtsam 1
28981 skämtsamheter 1
28982 skänka 3
28983 skänker 3
28984 skänkt 2
28985 skänkte 2
28986 skär 7
28987 skära 4
28988 skäras 3
28989 skärmen 6
28990 skärpa 7
28991 skärpas 2
28992 skärper 1
28993 skärpning 2
28994 skärpt 1
28995 skärpta 3
28996 skärrad 1
28997 skärs 3
28998 skärvor 1
28999 skådad 1
29000 skådade 1
29001 skådat 1
29002 skådespel 1
29003 skål 3
29004 skålade 1
29005 skålen 3
29006 skåp 2
29007 skåpdörr 1
29008 skåpet 3
29009 skåra 1
29010 sköldar 1
29011 sköldpaddan 1
29012 skölja 2
29013 sköljde 2
29014 sköna 1
29015 skönhet 6
29016 skönja 1
29017 skönjs 1
29018 skönt 1
29019 skör 1
29020 sköra 2
29021 skörd 3
29022 skörda 2
29023 skördar 1
29024 skördat 1
29025 skörden 2
29026 skörhet 1
29027 sköt 11
29028 sköta 14
29029 skötas 3
29030 sköter 4
29031 sköts 3
29032 skötsamma 1
29033 skötsel 2
29034 skötseln 1
29035 skötselnivå 1
29036 skött 3
29037 skötte 4
29038 skötts 2
29039 skövlade 1
29040 skövling 1
29041 skövlingen 1
29042 slag 45
29043 slagen 2
29044 slaget 8
29045 slagit 10
29046 slagkraftigt 1
29047 slagna 1
29048 slags 63
29049 slak 1
29050 slakt 3
29051 slaktar 2
29052 slaktarna 1
29053 slakten 1
29054 slaktprincip 1
29055 slaktprincipen 1
29056 slam 2
29057 slammer 2
29058 slampiga 1
29059 slamrade 1
29060 slamrande 1
29061 slamret 1
29062 slang 2
29063 slank 1
29064 slapp 1
29065 slappa 2
29066 slappare 1
29067 slapphet 5
29068 slappnade 1
29069 slarvig 1
29070 slarvigt 1
29071 slav 1
29072 slavar 2
29073 slaveri 2
29074 slem 1
29075 slemmet 1
29076 slemmiga 1
29077 slemtjockt 1
29078 slet 5
29079 slickade 2
29080 slingor 1
29081 slingrade 1
29082 slingrande 3
29083 slint 1
29084 slippa 9
29085 slipper 6
29086 slips 5
29087 slipsen 2
29088 slirar 1
29089 slita 2
29090 sliten 1
29091 sliter 2
29092 slits 1
29093 slitsammaste 1
29094 slockna 2
29095 slocknar 1
29096 slog 30
29097 slogan 1
29098 slogs 2
29099 slokande 1
29100 slopa 2
29101 slopandet 2
29102 slopar 1
29103 slopas 1
29104 slottspark 1
29105 slovenska 1
29106 slovensktalande 1
29107 slug 1
29108 slukade 1
29109 slukar 2
29110 slukas 1
29111 slumområden 1
29112 slump 7
29113 slumpat 1
29114 slumpen 2
29115 slumpmässig 1
29116 slumpmässiga 3
29117 slumpmässigt 1
29118 slumra 1
29119 slumrat 1
29120 slungades 1
29121 slunkit 1
29122 sluppit 1
29123 slussa 1
29124 slussas 1
29125 slut 82
29126 sluta 28
29127 slutade 1
29128 slutande 3
29129 slutandet 1
29130 slutanvändaren 1
29131 slutar 15
29132 slutare 1
29133 slutas 2
29134 slutat 5
29135 slutavtal 1
29136 slutdatum 3
29137 sluten 2
29138 slutenhet 1
29139 sluter 2
29140 slutet 82
29141 slutfasen 1
29142 slutför 1
29143 slutföra 6
29144 slutförande 1
29145 slutförandet 2
29146 slutföras 2
29147 slutförd 1
29148 slutfördes 1
29149 slutförs 2
29150 slutfört 4
29151 slutförts 4
29152 slutgiltig 2
29153 slutgiltiga 15
29154 slutgiltigt 8
29155 sluthanteringen 1
29156 slutit 6
29157 slutits 3
29158 slutkommentar 1
29159 slutkonsumenten 1
29160 slutlig 6
29161 slutliga 23
29162 slutligen 96
29163 slutligt 2
29164 slutmärke 3
29165 slutmärken 1
29166 slutmärkena 1
29167 slutmål 2
29168 slutmålet 1
29169 slutna 4
29170 slutomröstningen 3
29171 slutperioden 1
29172 slutpunkt 2
29173 slutresultat 1
29174 slutresultatet 3
29175 sluts 1
29176 slutsaten 1
29177 slutsats 12
29178 slutsatsen 19
29179 slutsatser 36
29180 slutsatserna 18
29181 slutstatusförhandlingarna 1
29182 sluttande 1
29183 sluttning 1
29184 sluttningarna 1
29185 sluttningen 4
29186 slutversionen 1
29187 slutändan 15
29188 slutänden 4
29189 slyngelstater 1
29190 släcka 3
29191 släcker 1
29192 släcks 1
29193 slädar 1
29194 släde 2
29195 släkt 1
29196 släkte 2
29197 släkten 1
29198 släktens 1
29199 släkting 1
29200 släktingar 4
29201 slänga 1
29202 slängde 6
29203 slänger 4
29204 slängs 2
29205 släp 1
29206 släpade 3
29207 släpades 1
29208 släpar 1
29209 släpets 1
29210 släppa 17
29211 släpper 5
29212 släpphänt 1
29213 släpphänta 1
29214 släpphänthet 1
29215 släpphäntheten 2
29216 släppområden 3
29217 släppområdets 1
29218 släpps 1
29219 släppt 2
29220 släppte 9
29221 släpptes 3
29222 släppts 1
29223 släta 3
29224 slätade 1
29225 slätnötta 1
29226 slätt 3
29227 slå 39
29228 slående 1
29229 slår 14
29230 slås 2
29231 slåss 3
29232 slösa 2
29233 slösade 1
29234 slösaktig 1
29235 slösar 1
29236 slösas 4
29237 slösat 1
29238 slösats 1
29239 slöseri 8
29240 slöseriet 1
29241 slöt 4
29242 slöts 1
29243 smak 1
29244 smakar 2
29245 smaken 1
29246 smaklösa 1
29247 smakämnen 1
29248 smal 6
29249 smala 2
29250 smalspårig 1
29251 smalt 1
29252 smart 4
29253 smarta 1
29254 smartare 1
29255 smekte 1
29256 smet 1
29257 smickrade 1
29258 smickrar 1
29259 smidesjärn 1
29260 smideskonstens 1
29261 smidig 2
29262 smidigare 1
29263 smidigt 1
29264 smids 1
29265 smita 1
29266 smitning 1
29267 smittad 4
29268 smittade 3
29269 smittades 1
29270 smittar 1
29271 smittas 1
29272 smittsam 2
29273 smittsamma 1
29274 smoking 1
29275 smokingjacka 1
29276 smuggelvaror 1
29277 smugglas 2
29278 smuggling 1
29279 smula 1
29280 smussla 1
29281 smusslande 1
29282 smuts 2
29283 smutsar 1
29284 smutsat 1
29285 smutsbruna 1
29286 smutsig 2
29287 smutsiga 5
29288 smutsigt 2
29289 smycka 1
29290 smycke 1
29291 smyg 1
29292 smyga 3
29293 smygande 1
29294 smyghandlare 1
29295 smäckra 1
29296 smädelse 1
29297 smädelser 1
29298 smäll 2
29299 smällde 1
29300 smält 1
29301 smälta 3
29302 smältande 1
29303 smältbar 1
29304 smärre 2
29305 smärta 7
29306 smärtar 1
29307 smärtas 1
29308 smärtfritt 1
29309 smärtsamma 1
29310 smärtsamt 4
29311 små 131
29312 små- 1
29313 småbarn 2
29314 småbrottslighet 1
29315 småfolket 1
29316 småföretag 8
29317 smågräl 1
29318 småhaiders 1
29319 småhuttra 1
29320 småjordbrukare 1
29321 småningom 14
29322 småpratade 1
29323 småpratar 1
29324 småsak 1
29325 småsaker 2
29326 småskaliga 2
29327 småskaligt 1
29328 småtrevligt 1
29329 smått 1
29330 smög 7
29331 smör 3
29332 smörgås 3
29333 smörgåsar 1
29334 smörgåspaket 1
29335 smörjan 1
29336 smörstekt 1
29337 snabb 19
29338 snabba 27
29339 snabbare 32
29340 snabbast 5
29341 snabbaste 3
29342 snabbhet 2
29343 snabbinsatscentral 1
29344 snabbinsatsstyrka 4
29345 snabbköp 1
29346 snabbt 155
29347 snabbvarningssystem 1
29348 snacka 1
29349 snake-heads 1
29350 snappa 1
29351 snar 10
29352 snarare 62
29353 snarast 30
29354 snaraste 1
29355 snarkade 1
29356 snarlika 1
29357 snart 78
29358 snaskiga 1
29359 snavande 1
29360 sned 1
29361 sneddade 1
29362 snedvrida 2
29363 snedvriden 2
29364 snedvrider 4
29365 snedvridning 12
29366 snedvridningar 6
29367 snedvridningarna 1
29368 snedvridningen 1
29369 snedvridningsriskerna 1
29370 snegla 1
29371 sneglade 1
29372 snett 5
29373 snickra 2
29374 snigeln 3
29375 snigelns 1
29376 snigelpost 1
29377 sniglar 1
29378 snikenhet 1
29379 snikenhetens 1
29380 snirkliga 1
29381 snobbig 1
29382 snoriga 1
29383 snort 1
29384 snubblade 1
29385 snubblande 1
29386 snuddar 1
29387 snurra 2
29388 snurrade 5
29389 snurrar 1
29390 snurrstolar 1
29391 snyftande 1
29392 snygg 3
29393 snyggt 2
29394 snäckdjuren 1
29395 snäll 5
29396 snälla 2
29397 snällt 1
29398 snärtar 1
29399 snäste 2
29400 snäv 1
29401 snävare 3
29402 snävt 1
29403 snåren 1
29404 snåriga 1
29405 snöiga 2
29406 snön 1
29407 snöret 2
29408 snörets 1
29409 snörpvad 2
29410 snörpvadfiske 1
29411 snövit 1
29412 snövitt 1
29413 so 1
29414 social 180
29415 social- 9
29416 sociala 401
29417 socialdemokrater 3
29418 socialdemokraterna 6
29419 socialdemokraternas 3
29420 socialdemokratin 1
29421 socialdemokratisk 3
29422 socialdemokratiska 30
29423 socialdemokratiske 1
29424 socialdemokratiskt 2
29425 socialdepartementet 1
29426 socialekonomisk 1
29427 socialekonomiska 2
29428 socialfonden 14
29429 socialfondens 3
29430 socialfrågor 15
29431 socialförsäkring 1
29432 socialförsäkringen 1
29433 socialförsäkringsfrågor 1
29434 socialförsäkringskostnaderna 1
29435 socialförsäkringsområdet 2
29436 socialförsäkringssystem 3
29437 socialförsäkringssystemen 3
29438 socialhjälp 1
29439 socialist 1
29440 socialister 8
29441 socialisterna 8
29442 socialisternas 1
29443 socialistgruppen 4
29444 socialistgruppens 1
29445 socialistisk 1
29446 socialistiska 19
29447 socialistkollegor 1
29448 socialistparti 1
29449 socialistpartiet 5
29450 socialistpartiets 2
29451 socialministrar 1
29452 socialpolitik 13
29453 socialpolitiken 17
29454 socialpolitikens 1
29455 socialpolitisk 1
29456 socialpolitiska 5
29457 socialrätt 1
29458 socialskyddet 2
29459 socialstatsmodellen 1
29460 socialstöd 3
29461 socialt 61
29462 socialtjänst 1
29463 society 3
29464 socio-ekonomiska 1
29465 socioekonomisk 1
29466 socioekonomiska 6
29467 sociokulturell 1
29468 sociologiska 1
29469 socker 1
29470 sockor 1
29471 sockrat 1
29472 sodomi 1
29473 soffa 1
29474 soffan 5
29475 soffbord 1
29476 soffbordet 2
29477 sofistikerade 2
29478 soft 1
29479 sola 2
29480 solblekta 1
29481 soldaten 1
29482 soldater 15
29483 soldaterna 2
29484 solen 10
29485 solens 1
29486 solfläck 1
29487 solglasögon 1
29488 solid 2
29489 solidarisera 1
29490 solidariserade 1
29491 solidarisk 8
29492 solidariska 4
29493 solidariskt 5
29494 solidaritet 62
29495 solidariteten 13
29496 solidaritetens 1
29497 solidaritetsarbetet 1
29498 solidaritetsförhållanden 1
29499 solidaritetssystem 1
29500 solidaritetsuttryck 1
29501 soliditet 1
29502 solig 3
29503 solkant 1
29504 solkungarnas 1
29505 solljus 1
29506 solljuset 4
29507 solnedgången 2
29508 solremsor 1
29509 solsken 4
29510 solskenet 3
29511 solstrålarna 1
29512 soluret 1
29513 som 11365
29514 somliga 13
29515 sommar 4
29516 sommaren 12
29517 sommarkvällarna 1
29518 sommarledighet 1
29519 sommarlov 2
29520 sommarlovet 1
29521 sommarnattens 1
29522 sommarsemester 1
29523 somnade 1
29524 son 14
29525 sonen 2
29526 sonens 1
29527 sons 1
29528 sopa 4
29529 sopade 1
29530 sopas 1
29531 sopats 1
29532 soppa 3
29533 soppan 1
29534 sopransångerskor 1
29535 soprantalare 1
29536 soptippen 1
29537 sorg 5
29538 sorger 1
29539 sorgfälligt 1
29540 sorgliga 2
29541 sorgligt 1
29542 sorgsen 1
29543 sorgsna 1
29544 sorlande 1
29545 sortens 10
29546 sorter 1
29547 sortera 4
29548 sortering 1
29549 sorters 2
29550 sorts 23
29551 sot 4
29552 sotet 1
29553 sov 4
29554 sova 4
29555 sovande 1
29556 sovit 1
29557 sovjetiska 2
29558 sovjettiden 1
29559 sovrum 1
29560 sovrummet 4
29561 sovrumsdörren 2
29562 sovvagn 1
29563 spanjor 6
29564 spanjorer 1
29565 spanjorerna 1
29566 spansk 4
29567 spanska 37
29568 spanske 1
29569 spanskt 2
29570 spara 18
29571 sparade 2
29572 sparande 4
29573 sparandet 1
29574 sparar 4
29575 sparare 1
29576 spararnas 2
29577 sparas 5
29578 sparat 1
29579 sparformer 1
29580 spark 1
29581 sparkade 1
29582 sparkar 2
29583 sparkas 1
29584 sparkassor 2
29585 sparmöjligheter 1
29586 sparpengar 2
29587 sparsamma 1
29588 sparvar 1
29589 special 4
29590 specialbestämmelser 4
29591 specialbilaga 1
29592 specialdomstolar 1
29593 specialeffekter 1
29594 specialfiske 1
29595 specialfordon 2
29596 specialförbanden 1
29597 specialinriktning 1
29598 specialiserad 2
29599 specialiserade 4
29600 specialiserat 2
29601 specialiseringen 1
29602 specialister 2
29603 specialistkompetens 1
29604 specialitet 1
29605 specialprogrammen 1
29606 specialtecken 1
29607 specialteckensekvenser 1
29608 specialutbildning 1
29609 speciell 17
29610 speciella 47
29611 speciellt 59
29612 specificera 3
29613 specificerade 1
29614 specificeranden 1
29615 specificerar 2
29616 specificeras 2
29617 specificering 2
29618 specifik 9
29619 specifika 50
29620 specifikation 2
29621 specifikationen 3
29622 specifikationer 1
29623 specifikt 16
29624 speditör 1
29625 speditörerna 1
29626 spegel 1
29627 spegeln 6
29628 spegla 1
29629 speglar 7
29630 speglas 1
29631 speglats 1
29632 spektakel 2
29633 spektakulär 2
29634 spektakulära 1
29635 spektrum 2
29636 spektrumet 3
29637 spekulation 1
29638 spekulationen 1
29639 spekulationer 1
29640 spekulationerna 1
29641 spekulativa 2
29642 spekulativt 1
29643 spekulera 2
29644 spekulerade 1
29645 spel 32
29646 spela 61
29647 spelad 1
29648 spelade 10
29649 spelar 43
29650 spelare 1
29651 spelas 1
29652 spelat 13
29653 spelbrickor 1
29654 spelen 2
29655 spelet 4
29656 spelfält 1
29657 spelfältet 1
29658 spelkort 1
29659 spelpjäser 1
29660 spelplan 1
29661 spelregler 8
29662 spelreglerna 2
29663 spelrum 1
29664 spelrummet 1
29665 spendera 3
29666 spenderar 3
29667 spenderas 2
29668 spets 1
29669 spetsade 1
29670 spetsen 6
29671 spetsföretag 1
29672 spetsig 1
29673 spetsiga 3
29674 spettet 1
29675 spika 1
29676 spilla 1
29677 spillo 2
29678 spillolja 2
29679 spillror 1
29680 spills 2
29681 spindelnätet 1
29682 spindlar 1
29683 spionerade 1
29684 spiral 2
29685 spiror 1
29686 spis 1
29687 spisar 1
29688 spisarna 1
29689 spiselhyllan 2
29690 spisen 1
29691 spjut 2
29692 spjutspets 1
29693 splay 1
29694 split 2
29695 splitterny 1
29696 splittra 1
29697 splittrad 3
29698 splittrade 3
29699 splittras 4
29700 splittrat 2
29701 splittrats 1
29702 splittring 5
29703 spola 1
29704 spolas 3
29705 spongiform 1
29706 sponsorer 1
29707 sponsrad 1
29708 spontan 2
29709 spontana 1
29710 spontaniteten 1
29711 spontant 4
29712 sporadisk 1
29713 sporra 1
29714 sporre 2
29715 sporren 1
29716 sport 2
29717 sporta 1
29718 sportavsnittet 1
29719 sportbåtar 1
29720 sportfantaster 1
29721 sportfiskare 1
29722 spots 1
29723 sprack 3
29724 sprakade 1
29725 sprang 10
29726 spratt 1
29727 spred 4
29728 spreds 4
29729 spreta 1
29730 spricka 3
29731 sprickan 2
29732 spricker 1
29733 sprickor 1
29734 sprida 9
29735 spridande 1
29736 spridandet 1
29737 spridas 7
29738 spridd 1
29739 spridda 1
29740 sprider 12
29741 spridits 2
29742 spridning 17
29743 spridningen 5
29744 spridningsreglerna 1
29745 sprids 7
29746 springa 6
29747 springande 3
29748 springares 1
29749 springpojke 1
29750 sprit 2
29751 spritts 1
29752 sprudlar 1
29753 sprungen 1
29754 sprungit 1
29755 sprutade 1
29756 sprutas 1
29757 sprutt 1
29758 spräcka 1
29759 spräckt 1
29760 spräckte 1
29761 sprängande 1
29762 sprängämnen 1
29763 språk 31
29764 språkbruk 3
29765 språken 1
29766 språket 8
29767 språkets 1
29768 språkgrupper 1
29769 språklig 3
29770 språkliga 3
29771 språkområden 1
29772 språkområdena 1
29773 språkversioner 1
29774 språng 2
29775 spröd 1
29776 spurt 1
29777 spurts 1
29778 spy 2
29779 spädbarn 1
29780 spädbarns 2
29781 spädbarnsdödligheten 1
29782 spänd 3
29783 spända 2
29784 spände 2
29785 spänna 2
29786 spännande 11
29787 spänner 1
29788 spänning 9
29789 spänningar 7
29790 spänningarna 3
29791 spänningen 1
29792 spänningsfält 1
29793 spänningsförhållandet 1
29794 spänst 1
29795 spänt 2
29796 spär 1
29797 spärr 1
29798 spärrad 1
29799 spärrar 2
29800 spärras 1
29801 spärreld 1
29802 spådomar 1
29803 spår 11
29804 spåra 4
29805 spåras 1
29806 spårbarhet 4
29807 spåren 1
29808 spåret 1
29809 spårning 1
29810 spöke 3
29811 spöken 1
29812 spöklika 1
29813 spökstäder 1
29814 spörsmålet 1
29815 srilankesiska 1
29816 stab 2
29817 stabil 9
29818 stabila 6
29819 stabilare 1
29820 stabilisera 3
29821 stabiliserande 1
29822 stabiliseras 1
29823 stabilisering 4
29824 stabiliseringen 1
29825 stabiliserings- 14
29826 stabiliseringspakten 1
29827 stabiliseringsprocess 1
29828 stabiliseringssträvan 1
29829 stabilitet 38
29830 stabiliteten 15
29831 stabilitetsfaktor 1
29832 stabilitetskursen 1
29833 stabilitetslänk 1
29834 stabilitetspakt 4
29835 stabilitetspakten 20
29836 stabilitetsplanen 1
29837 stabilitetspolitik 1
29838 stabilitetspolitiken 2
29839 stabilt 5
29840 stablitetskultur 1
29841 stack 3
29842 stackars 5
29843 stackatokaskader 1
29844 stad 17
29845 staden 18
29846 stadens 1
29847 stadga 40
29848 stadgan 41
29849 stadgans 1
29850 stadgar 4
29851 stadgehänseende 1
29852 stadier 1
29853 stadiet 3
29854 stadig 2
29855 stadigt 5
29856 stadigvarande 1
29857 stadion 1
29858 stadium 8
29859 stads 1
29860 stads- 2
29861 stadsbefolkningen 1
29862 stadsboende 1
29863 stadsbor 1
29864 stadscentrum 1
29865 stadsdel 1
29866 stadsdelar 2
29867 stadsdelarna 2
29868 stadsdelen 1
29869 stadsförnyelse 1
29870 stadskärnor 2
29871 stadsmiljö 2
29872 stadsmiljögrupp 1
29873 stadsmiljöinitiativ 1
29874 stadsmiljöinitiativet 2
29875 stadsmiljön 1
29876 stadsområde 3
29877 stadsområden 12
29878 stadsområdena 3
29879 stadsområdet 1
29880 stadsplaneringen 1
29881 stadspolitik 1
29882 stadspolitiken 1
29883 stadsrelaterade 1
29884 stadsutveckling 3
29885 stagnation 2
29886 stagnerar 1
29887 stagnerat 2
29888 staka 1
29889 stakeholder 1
29890 stakeholders 1
29891 stalinistiska 1
29892 stalinistiskt 1
29893 stalldörren 1
29894 stammarna 1
29895 stammen 3
29896 stampa 1
29897 stampande 1
29898 stampar 1
29899 stan 7
29900 standard 18
29901 standardanpassningen 1
29902 standardbaserat 1
29903 standarden 2
29904 standarder 8
29905 standardernas 1
29906 standardfilformat 1
29907 standardformatmall 1
29908 standardformuleringar 1
29909 standardfrågeläget 1
29910 standardhöjande 1
29911 standardinstallationen 1
29912 standardinställning 1
29913 standardinställningen 1
29914 standardiserade 4
29915 standardiseras 1
29916 standardisering 3
29917 standardiseringar 2
29918 standardiseringen 1
29919 standardiseringskommittén 3
29920 standardiseringssträvandena 2
29921 standardkontot 1
29922 standards 1
29923 standardspråket 2
29924 stanken 1
29925 stanna 19
29926 stannade 12
29927 stannande 1
29928 stannar 7
29929 stannat 6
29930 stans 1
29931 staplade 1
29932 staplades 1
29933 stark 44
29934 starka 40
29935 starkare 24
29936 starkast 4
29937 starkaste 5
29938 starke 2
29939 starkt 76
29940 starmade 1
29941 stars 1
29942 start 2
29943 start- 2
29944 start-up-fenomenet 1
29945 start-up-företags 1
29946 starta 17
29947 startade 4
29948 startades 2
29949 startar 4
29950 startas 3
29951 startat 3
29952 startats 3
29953 starten 5
29954 startkapital 1
29955 startmärke 2
29956 startplatta 1
29957 startpunkten 2
29958 stass 1
29959 stat 44
29960 staten 38
29961 statens 9
29962 stater 56
29963 stater-nationer 1
29964 staterna 104
29965 staternas 31
29966 staters 2
29967 station 2
29968 stationen 14
29969 stationens 3
29970 stationerade 1
29971 stationerna 1
29972 stationsvagn 1
29973 stationära 1
29974 statister 1
29975 statistik 14
29976 statistiken 2
29977 statistikens 1
29978 statistisk 3
29979 statistiska 7
29980 statistiskt 4
29981 statlig 12
29982 statliga 75
29983 statligt 28
29984 stats 4
29985 stats- 10
29986 statsbal 1
29987 statsbalen 1
29988 statsbudgeten 1
29989 statschefen 1
29990 statschefer 2
29991 statschefers 1
29992 statsfinanser 1
29993 statsförbund 1
29994 statsgrundandet 1
29995 statskapitalism 1
29996 statskassan 2
29997 statskuppen 1
29998 statslösa 1
29999 statsmakt 6
30000 statsmakten 2
30001 statsmaktens 1
30002 statsmakterna 2
30003 statsminister 1
30004 statsministern 1
30005 statsministrarnas 1
30006 statsmonopolet 1
30007 statsmonopolets 1
30008 statsobligationer 1
30009 statssekreteraren 1
30010 statssekreterarens 1
30011 statsskulden 1
30012 statsskulder 1
30013 statsstöd 10
30014 statsstöden 4
30015 statsstödens 3
30016 statsstödet 1
30017 statsstödspolitiken 1
30018 statssäkerheten 1
30019 statstelevision 1
30020 statstjänstemän 1
30021 statsutgifter 1
30022 statsvetare 1
30023 statsvetenskapens 1
30024 statsåklagaren 1
30025 statsöverhuvudena 1
30026 statuera 2
30027 statuerar 1
30028 status 15
30029 statusen 2
30030 stavar 2
30031 stavningsarbete 1
30032 stearinljus 2
30033 steering 1
30034 steg 132
30035 stegade 1
30036 stegen 8
30037 steget 9
30038 stegrades 1
30039 stegsumman 1
30040 stegvis 1
30041 stek 1
30042 stekflott 1
30043 stekhus 1
30044 stekpannan 2
30045 stel 4
30046 stela 5
30047 stella 2
30048 stelt 3
30049 sten 9
30050 stenar 2
30051 stenbeläggning 1
30052 stenbrott 1
30053 stenbyggnader 1
30054 stendövt 1
30055 stenen 1
30056 stenfasaden 1
30057 stenhårda 1
30058 steniga 1
30059 stenigt 1
30060 stenkall 1
30061 stenkolen 1
30062 stenkolsindustrierna 1
30063 stenkolsindustrin 2
30064 stenmur 1
30065 stenplattor 1
30066 stereotypa 1
30067 stereotyper 2
30068 steril 1
30069 stetoskopet 1
30070 stick 3
30071 sticka 6
30072 stickade 1
30073 stickande 1
30074 stickare 1
30075 sticker 3
30076 sticket 2
30077 stickord 1
30078 stickprovskontroll 1
30079 stickprovskontroller 1
30080 stickprovstest 1
30081 stickprovsundersökningar 1
30082 stifta 3
30083 stiftar 1
30084 stig 2
30085 stiga 5
30086 stigande 3
30087 stigar 2
30088 stigen 2
30089 stiger 5
30090 stigit 10
30091 stigmatiserat 1
30092 stil 5
30093 stilen 1
30094 stilig 2
30095 stiliserade 1
30096 stilla 9
30097 stillasittande 1
30098 stillastående 2
30099 stillhet 3
30100 stillheten 1
30101 stillsamt 2
30102 stilmall 1
30103 stilmallen 1
30104 stimulans 8
30105 stimulansen 3
30106 stimulanser 3
30107 stimulansåtgärder 2
30108 stimulansåtgärderna 1
30109 stimulera 13
30110 stimulerande 7
30111 stimulerar 3
30112 stimulerat 1
30113 stimulering 1
30114 stinkande 1
30115 stinker 1
30116 stint 1
30117 stipulerade 1
30118 stirra 1
30119 stirrade 11
30120 stirrande 1
30121 stirrar 2
30122 stirrat 1
30123 stjäl 1
30124 stjäla 2
30125 stjärna 2
30126 stjärnfisk 1
30127 stjärnor 3
30128 stjärnorna 3
30129 stjärnornas 1
30130 stjärt 1
30131 stjärten 1
30132 stockflottorna 1
30133 stockning 1
30134 stocks 1
30135 stod 61
30136 stoft 1
30137 stoftblandning 1
30138 stoftkorn 1
30139 stol 2
30140 stolar 3
30141 stolarna 1
30142 stolen 6
30143 stolsitsen 1
30144 stolt 15
30145 stolta 5
30146 stolte 1
30147 stolthet 10
30148 stoltsera 2
30149 stoltserar 1
30150 stopp 29
30151 stoppa 12
30152 stoppade 3
30153 stoppades 2
30154 stoppar 1
30155 stoppas 9
30156 stoppat 1
30157 stoppats 1
30158 stor 324
30159 stora 355
30160 storartad 1
30161 storartat 3
30162 stordrifts- 1
30163 stordriftsfördelar 1
30164 stordriftsfördelarna 1
30165 store 1
30166 storföretag 2
30167 storföretagens 1
30168 storhet 2
30169 storheter 1
30170 storhetsvansinne 1
30171 storkapitalet 1
30172 storkapitalets 2
30173 storkonsument 1
30174 storlek 10
30175 storlekar 1
30176 storleken 5
30177 storleksordningen 3
30178 storleksskaften 1
30179 storm 2
30180 storma 1
30181 stormakt 1
30182 stormakterna 1
30183 stormar 8
30184 stormarknader 2
30185 stormarna 12
30186 stormarnas 1
30187 stormen 6
30188 stormens 1
30189 stormfloden 1
30190 stormfällda 1
30191 stormvind 1
30192 storsinta 1
30193 storskalig 1
30194 storskaliga 4
30195 storskalighet 1
30196 storslaget 1
30197 storslagna 2
30198 storstadsförorter 1
30199 storstäderna 3
30200 stort 135
30201 stortårna 1
30202 storvulen 1
30203 story 1
30204 straff 10
30205 straff- 2
30206 straffa 5
30207 straffas 4
30208 straffats 1
30209 straffbar 2
30210 straffbara 1
30211 straffbarheten 1
30212 straffbart 1
30213 straffbestämmelser 1
30214 straffet 2
30215 strafflagstiftning 2
30216 straffläger 1
30217 strafflöshet 1
30218 straffprocessrätten 1
30219 straffprocessrättsligt 1
30220 straffrihet 1
30221 straffriheten 1
30222 straffrätt 10
30223 straffrätten 12
30224 straffrättens 3
30225 straffrättslig 3
30226 straffrättsliga 32
30227 straffrättsligt 10
30228 straffrättsområdet 1
30229 stragglande 1
30230 stram 3
30231 strama 2
30232 stramhet 1
30233 strand 1
30234 stranda 1
30235 stranden 4
30236 strandremsa 4
30237 strandremsan 2
30238 strandremsans 1
30239 strategi 88
30240 strategidokument 2
30241 strategier 37
30242 strategierna 3
30243 strategin 19
30244 strategiplanering 1
30245 strategisk 11
30246 strategiska 51
30247 strategiskt 13
30248 strax 13
30249 streck 1
30250 strecksats 1
30251 stress 1
30252 stretar 1
30253 stretch 1
30254 strid 24
30255 strida 6
30256 stridande 1
30257 striden 3
30258 strider 25
30259 stridigheten 1
30260 stridslystet 1
30261 stridsropet 1
30262 stridsvagnar 1
30263 strikt 25
30264 strikta 17
30265 striktare 6
30266 strimma 2
30267 strimman 1
30268 strimmorna 1
30269 stringens 1
30270 stringentare 1
30271 stripes 1
30272 stripigt 1
30273 strukits 2
30274 struktur 34
30275 strukturanpassningen 1
30276 strukturell 7
30277 strukturella 25
30278 strukturellt 6
30279 strukturen 19
30280 strukturer 37
30281 strukturera 2
30282 strukturerad 3
30283 strukturerande 2
30284 strukturerar 1
30285 struktureras 2
30286 strukturerat 6
30287 struktureringen 1
30288 strukturerna 8
30289 strukturers 1
30290 strukturfonden 3
30291 strukturfonder 18
30292 strukturfonderna 96
30293 strukturfonderna- 1
30294 strukturfondernas 6
30295 strukturfondsförordningen 1
30296 strukturfondsmedel 1
30297 strukturfondsprogram 1
30298 strukturfondsprogrammen 2
30299 strukturfondsrunda 1
30300 strukturfondsstödet 1
30301 strukturformerna 2
30302 strukturförändringen 1
30303 strukturmässig 1
30304 strukturpolitik 8
30305 strukturpolitiken 5
30306 strukturprojekt 1
30307 strukturreformer 3
30308 strukturstramhet 1
30309 strukturstöd 4
30310 strukturstöden 1
30311 strukturutgifterna 1
30312 strukturutveckling 2
30313 strukturåtgärderna 1
30314 strumpor 4
30315 strumporna 1
30316 strumpstickor 1
30317 strumpsömmar 1
30318 strunt 1
30319 strunta 5
30320 struntar 3
30321 struntat 1
30322 struntprat 3
30323 strupen 1
30324 struts 1
30325 stryk 1
30326 stryka 5
30327 strykas 2
30328 strykningen 1
30329 stryks 3
30330 stryps 1
30331 strypt 1
30332 sträck 1
30333 sträcka 9
30334 sträckan 1
30335 sträcker 9
30336 sträckor 1
30337 sträckte 6
30338 stränder 10
30339 stränderna 6
30340 sträng 8
30341 stränga 15
30342 strängare 5
30343 strängaste 2
30344 stränghet 4
30345 strängt 9
30346 sträva 16
30347 strävade 2
30348 strävan 27
30349 strävanden 7
30350 strävandena 1
30351 strävar 20
30352 strävat 1
30353 strået 2
30354 strålade 1
30355 strålande 2
30356 strålar 1
30357 stråle 1
30358 strålkastare 1
30359 strålkastaren 1
30360 strålkastarljuset 1
30361 strålning 1
30362 strålskydd 1
30363 strödde 1
30364 strök 1
30365 ströks 1
30366 ström 7
30367 strömmade 3
30368 strömmande 2
30369 strömmarna 1
30370 strömningar 4
30371 strömningarna 1
30372 strömningen 2
30373 ströva 1
30374 strövade 1
30375 stuckit 1
30376 student 3
30377 studenten 1
30378 studenter 3
30379 studenterna 1
30380 studentskan 1
30381 studera 2
30382 studerade 3
30383 studerar 4
30384 studeras 2
30385 studerat 3
30386 studie 6
30387 studiebesök 1
30388 studiedag 1
30389 studien 1
30390 studieprogram 1
30391 studier 17
30392 studsade 2
30393 stugor 1
30394 stum 3
30395 stumme 1
30396 stund 32
30397 stundande 3
30398 stunden 3
30399 stunder 4
30400 stunderna 1
30401 stundtals 1
30402 stuvade 1
30403 stycke 4
30404 stycken 3
30405 styckena 2
30406 stycket 4
30407 stympad 2
30408 stympningen 1
30409 styr 6
30410 styra 19
30411 styrande 2
30412 styras 6
30413 styrd 1
30414 styrda 1
30415 styrde 4
30416 styre 3
30417 styrekonomen 3
30418 styrelse 3
30419 styrelsebeslut 1
30420 styrelseformer 1
30421 styrelseformerna 1
30422 styrelsen 3
30423 styrelser 1
30424 styrelseskick 1
30425 styret 2
30426 styrets 1
30427 styrka 13
30428 styrkan 4
30429 styrkeförhållandena 2
30430 styrkeposition 1
30431 styrketest 1
30432 styrkommittéerna 1
30433 styrkor 15
30434 styrkorna 5
30435 styrning 2
30436 styrningen 2
30437 styrs 6
30438 styrt 3
30439 styva 1
30440 styvsint 1
30441 styvt 1
30442 städ 1
30443 städa 5
30444 städade 2
30445 städat 2
30446 städer 29
30447 städerna 29
30448 städernas 5
30449 städers 2
30450 städning 1
30451 ställ 1
30452 ställa 99
30453 ställas 32
30454 ställda 2
30455 ställde 28
30456 ställdes 6
30457 ställe 16
30458 ställen 9
30459 ställer 69
30460 stället 139
30461 ställning 73
30462 ställningar 1
30463 ställningen 1
30464 ställningstagande 12
30465 ställningstaganden 4
30466 ställningstagandet 1
30467 ställs 30
30468 ställt 24
30469 ställts 8
30470 stämde 3
30471 stämma 6
30472 stämmer 35
30473 stämning 1
30474 stämningen 3
30475 stämningsansökningar 1
30476 stämpling 1
30477 ständig 7
30478 ständiga 15
30479 ständigt 45
30480 stänga 3
30481 stängda 3
30482 stängde 5
30483 stängdes 1
30484 stänger 3
30485 stängerna 1
30486 stängning 3
30487 stängningen 2
30488 stängs 3
30489 stängsel 1
30490 stängts 3
30491 stänkte 2
30492 stärka 65
30493 stärkande 6
30494 stärkandet 4
30495 stärkas 8
30496 stärkelsevit 1
30497 stärker 9
30498 stärks 5
30499 stärkt 3
30500 stärkts 2
30501 stäv 3
30502 stävja 1
30503 stävjas 1
30504 stå 68
30505 stående 7
30506 stål 1
30507 stålföretag 5
30508 stålgemenskapen 1
30509 stålindustrin 23
30510 stålindustrins 2
30511 stålsektorn 4
30512 stålverk 2
30513 stålverket 2
30514 stålverksanläggningar 1
30515 stånd 61
30516 ståndpunkt 139
30517 ståndpunkten 65
30518 ståndpunkter 41
30519 ståndpunkterna 5
30520 ståndpunktstagande 1
30521 stång 1
30522 står 258
30523 ståtlig 2
30524 stått 18
30525 stöd 348
30526 stöd- 1
30527 stödbehov 1
30528 stödberättigade 7
30529 stödberättigande 1
30530 stödd 3
30531 stödda 1
30532 stödde 6
30533 stöddes 1
30534 stöden 26
30535 stöder 166
30536 stödet 51
30537 stödets 1
30538 stödformer 1
30539 stödinstrument 1
30540 stödja 167
30541 stödjande 3
30542 stödjas 14
30543 stödjer 5
30544 stödkategorier 1
30545 stödköper 1
30546 stödmedlen 1
30547 stödmekanismer 1
30548 stödmottagaren 1
30549 stödmöjligheter 1
30550 stödnivån 2
30551 stödområden 1
30552 stödområdena 1
30553 stödpolitik 1
30554 stödprogram 5
30555 stödpunkt 1
30556 stödpunkten 1
30557 stödram 1
30558 stödramar 1
30559 stöds 16
30560 stödsystem 3
30561 stödsystemet 1
30562 stödsänkningarna 1
30563 stödverktygen 1
30564 stödyta 1
30565 stödåtgärder 11
30566 stödåtgärderna 2
30567 stöld 3
30568 stönade 1
30569 stönande 1
30570 stöpa 2
30571 stöpsleven 1
30572 stör 6
30573 störa 3
30574 störande 3
30575 störas 1
30576 störd 2
30577 störde 3
30578 störning 1
30579 störningar 5
30580 störningarna 1
30581 större 209
30582 störs 2
30583 störst 9
30584 största 106
30585 störste 1
30586 störta 3
30587 störtade 2
30588 störtflod 1
30589 stöt 3
30590 stöta 2
30591 stötande 1
30592 stöten 1
30593 stöter 2
30594 stötestenarna 1
30595 stötfångare 1
30596 stött 19
30597 stötta 2
30598 stöttat 2
30599 stötte 5
30600 stöttepelare 1
30601 stöttepelaren 1
30602 stötts 2
30603 stövlar 1
30604 sua 1
30605 sub 1
30606 subject 1
30607 subjekt 1
30608 subjektiva 1
30609 sublima 1
30610 subsidaritetsprincipen 2
30611 subsidiaritet 10
30612 subsidiariteten 11
30613 subsidiaritets- 1
30614 subsidiaritetsaltaret 1
30615 subsidiaritetsfrågor 2
30616 subsidiaritetsprincip 1
30617 subsidiaritetsprincipen 28
30618 subsidiaritetsprinciper 1
30619 subsidiär 1
30620 substans 2
30621 substansen 1
30622 substantiella 2
30623 substantiellt 1
30624 substitut 2
30625 subtila 1
30626 subvention 1
30627 subventioner 12
30628 subventionera 3
30629 subventionerade 1
30630 subventionerar 1
30631 subventioneras 1
30632 subventionerna 2
30633 subventionskonkurrens 1
30634 successiv 2
30635 successiva 4
30636 successivt 7
30637 sucka 1
30638 suckade 3
30639 suckades 1
30640 suckar 1
30641 sudaneserna 1
30642 sudda 2
30643 suddades 1
30644 suddig 1
30645 suger 1
30646 sugs 1
30647 summa 6
30648 summan 2
30649 summarisk 1
30650 summera 1
30651 summertonen 1
30652 summor 13
30653 sund 4
30654 sunda 7
30655 sundare 3
30656 sundaste 1
30657 sundhet 1
30658 sunt 4
30659 supa 1
30660 superdistinguished 1
30661 supereuropéerna 1
30662 supermakt 2
30663 superstat 1
30664 supranationell 1
30665 surrad 1
30666 surrade 3
30667 surrande 1
30668 surrogat 1
30669 surrogatfader 2
30670 surögt 1
30671 susade 1
30672 suspekta 1
30673 suspenderas 1
30674 suspensiv 1
30675 suttit 7
30676 suverän 2
30677 suveräna 5
30678 suveränitet 19
30679 suveräniteten 6
30680 suveränt 1
30681 svag 11
30682 svaga 12
30683 svagare 10
30684 svagares 1
30685 svagaste 6
30686 svaghet 12
30687 svagheten 3
30688 svagheter 4
30689 svagheterna 3
30690 svagt 4
30691 svaj 1
30692 svajade 1
30693 sval 1
30694 svala 1
30695 svalde 1
30696 svalka 1
30697 svansar 1
30698 svansen 2
30699 svar 121
30700 svara 45
30701 svarade 24
30702 svarande 1
30703 svarar 18
30704 svarat 8
30705 svaren 8
30706 svaret 25
30707 svaromål 1
30708 svars 9
30709 svarstider 1
30710 svarston 1
30711 svart 21
30712 svarta 26
30713 svartas 1
30714 svarte 1
30715 svartingar 2
30716 svartingarna 1
30717 svartjobb 1
30718 svartklädda 2
30719 svartkonst 1
30720 svartkonstnären 1
30721 svartlista 1
30722 svartröd 1
30723 svartsjuka 1
30724 svassa 1
30725 svavelhalt 1
30726 svavelhalten 1
30727 svek 3
30728 svekfullt 1
30729 svensk 4
30730 svenska 22
30731 svenskarna 1
30732 svenske 1
30733 svensken 1
30734 svenskt 1
30735 svepande 1
30736 svepskäl 2
30737 svepte 6
30738 svett 3
30739 svetten 2
30740 svettglänsande 1
30741 svikit 1
30742 svinaktigt 1
30743 svindel 2
30744 svindlande 1
30745 svinstia 1
30746 svischade 1
30747 sviterna 1
30748 svurit 1
30749 svälja 1
30750 svällande 1
30751 svält 5
30752 svälta 1
30753 svältsituationer 1
30754 svämmade 1
30755 svämmar 1
30756 svänga 1
30757 svängande 2
30758 svängd 1
30759 svängde 4
30760 svängningar 1
30761 svängrum 1
30762 svär 1
30763 svärd 2
30764 svärdet 1
30765 svärta 2
30766 svärtas 1
30767 sväva 1
30768 svävade 3
30769 svävande 4
30770 svåger 1
30771 svågerpolitik 3
30772 svål 1
30773 svångrems- 1
30774 svår 28
30775 svåra 45
30776 svårare 11
30777 svårartade 1
30778 svåraste 2
30779 svårbedömbara 1
30780 svårbegriplig 2
30781 svårhanterliga 1
30782 svårighet 2
30783 svårigheten 5
30784 svårigheter 70
30785 svårigheterna 13
30786 svårligen 1
30787 svårlöst 1
30788 svårlösta 1
30789 svårmod 1
30790 svårt 105
30791 svårtolkat 1
30792 svåröverskådligt 1
30793 svåröverstigliga 1
30794 syd 1
30795 sydafrikanen 2
30796 sydafrikanens 1
30797 sydafrikanerna 1
30798 sydafrikanska 1
30799 sydamerikanska 1
30800 sydeuropeiska 1
30801 sydkusten 1
30802 sydlig 1
30803 sydliga 2
30804 sydligt 1
30805 sydvästra 2
30806 sydöstra 10
30807 syfta 2
30808 syftade 5
30809 syftande 1
30810 syftar 79
30811 syfte 85
30812 syften 13
30813 syftena 2
30814 syftet 41
30815 sykomorträ 1
30816 symbol 8
30817 symbolen 1
30818 symboler 1
30819 symbolerna 1
30820 symbolisera 1
30821 symboliserar 1
30822 symbolisk 5
30823 symboliska 4
30824 symboliskt 1
30825 symbolism 1
30826 symfoniorkestrar 1
30827 sympati 10
30828 sympatier 1
30829 sympatiserade 1
30830 sympatiserar 3
30831 sympatiskt 2
30832 sympatiyttring 1
30833 symptom 3
30834 symptomatiska 1
30835 symptomen 1
30836 symtom 2
30837 syn 32
30838 syna 1
30839 synar 1
30840 synas 3
30841 synd 13
30842 syndabock 1
30843 syndabockar 2
30844 syndar 1
30845 synder 1
30846 syndikalister 2
30847 syndromet 1
30848 synen 4
30849 synergi 1
30850 synergieffekter 3
30851 synergierna 1
30852 synergism 1
30853 synes 4
30854 synfält 1
30855 synhåll 2
30856 synkronicitet 1
30857 synkroniserad 1
30858 synkroniseringen 1
30859 synlig 5
30860 synliga 7
30861 synligare 1
30862 synligaste 1
30863 synliggörs 1
30864 synligt 2
30865 synnerhet 163
30866 synnerligen 17
30867 synonym 1
30868 synonymt 1
30869 synpunkt 18
30870 synpunkten 7
30871 synpunkter 47
30872 synpunkterna 2
30873 syns 2
30874 synsätt 13
30875 synsättet 1
30876 syntax-regler 1
30877 syntes 5
30878 syntetiska 1
30879 synvinkel 26
30880 synvinkeln 8
30881 synvinklar 1
30882 syrier 1
30883 syrierna 3
30884 syriska 4
30885 syriske 1
30886 sysselsatt 4
30887 sysselsatta 3
30888 sysselsätta 2
30889 sysselsätter 4
30890 sysselsättning 195
30891 sysselsättningen 87
30892 sysselsättningens 3
30893 sysselsättnings- 3
30894 sysselsättningsargumentet 1
30895 sysselsättningsbas 1
30896 sysselsättningsdrivande 1
30897 sysselsättningsfaktor 1
30898 sysselsättningsfluktuationerna 1
30899 sysselsättningsfrämjande 2
30900 sysselsättningsfrågan 2
30901 sysselsättningsförhållanden 1
30902 sysselsättningsförmåga 3
30903 sysselsättningsgrad 4
30904 sysselsättningsinitiativ 1
30905 sysselsättningsinitiativen 1
30906 sysselsättningskvaliteten 1
30907 sysselsättningsläget 1
30908 sysselsättningsmodeller 1
30909 sysselsättningsmöjligheter 2
30910 sysselsättningsnivå 4
30911 sysselsättningsnivåer 1
30912 sysselsättningsnivåerna 1
30913 sysselsättningsnivån 4
30914 sysselsättningsområden 1
30915 sysselsättningsområdet 2
30916 sysselsättningspaketet 1
30917 sysselsättningspakten 1
30918 sysselsättningspakterna 1
30919 sysselsättningsplaner 1
30920 sysselsättningspolitik 11
30921 sysselsättningspolitiken 15
30922 sysselsättningspolitiska 6
30923 sysselsättningspotential 2
30924 sysselsättningsproblem 2
30925 sysselsättningsproblematiken 2
30926 sysselsättningsprogrammen 1
30927 sysselsättningsrapporten 2
30928 sysselsättningssamarbetet 1
30929 sysselsättningsskapande 6
30930 sysselsättningsskydd 1
30931 sysselsättningsstrategi 2
30932 sysselsättningsstrategier 1
30933 sysselsättningsstrategin 7
30934 sysselsättningsstrategins 1
30935 sysselsättningstoppmötet 1
30936 sysselsättningsvänliga 1
30937 sysselsättningsåtgärder 1
30938 sysselsättningsåtgärderna 1
30939 sysselsättningsökningen 1
30940 syssla 3
30941 sysslade 3
30942 sysslar 9
30943 sysslolösa 3
30944 system 175
30945 systemadministratör 1
30946 systemadministratören 1
30947 systematisera 1
30948 systematisk 10
30949 systematiska 2
30950 systematiskt 12
30951 systemen 20
30952 systemet 80
30953 systemets 1
30954 systemmodernisering 1
30955 systemutveckling 1
30956 systemändring 2
30957 systemändringen 1
30958 syster 3
30959 systerfartyg 1
30960 systern 1
30961 systerskap 1
30962 systerson 1
30963 systrar 5
30964 säden 1
30965 sädesbåtarna 1
30966 säg 4
30967 säga 539
30968 sägas 12
30969 säger 249
30970 sägs 17
30971 säker 73
30972 säkerhet 144
30973 säkerheten 48
30974 säkerhetens 2
30975 säkerhets 2
30976 säkerhets- 8
30977 säkerhetsanordning 1
30978 säkerhetsargument 1
30979 säkerhetsaspekten 1
30980 säkerhetsbestämmelser 2
30981 säkerhetsbestämmelserna 1
30982 säkerhetsbältet 1
30983 säkerhetsfrågan 2
30984 säkerhetsfrågor 2
30985 säkerhetsfångar 1
30986 säkerhetsföreskrifterna 1
30987 säkerhetsförhållandena 1
30988 säkerhetsgarantierna 2
30989 säkerhetsgränsen 1
30990 säkerhetshänsyn 1
30991 säkerhetsinsatserna 1
30992 säkerhetsinställningar 1
30993 säkerhetsintresse 1
30994 säkerhetskontrollerna 1
30995 säkerhetskopia 1
30996 säkerhetskopian 1
30997 säkerhetskrav 1
30998 säkerhetskriser 1
30999 säkerhetsläget 2
31000 säkerhetsnivå 1
31001 säkerhetsnivån 1
31002 säkerhetsnormer 2
31003 säkerhetsnätet 1
31004 säkerhetsorganisation 1
31005 säkerhetspolitik 15
31006 säkerhetspolitiken 9
31007 säkerhetspolitikens 1
31008 säkerhetspolitisk 1
31009 säkerhetsproblem 2
31010 säkerhetsproblemen 1
31011 säkerhetsrisk 3
31012 säkerhetsrisker 1
31013 säkerhetsråd 7
31014 säkerhetsrådet 2
31015 säkerhetsrådets 4
31016 säkerhetsrådgivare 12
31017 säkerhetsrådgivarna 1
31018 säkerhetsråds 1
31019 säkerhetsskäl 1
31020 säkerhetsstyrka 1
31021 säkerhetsstyrkans 1
31022 säkerhetsställande 1
31023 säkerhetssystemet 1
31024 säkerhetstjänst 1
31025 säkerhetsventil 1
31026 säkerhetsåtgärd 1
31027 säkerhetsåtgärderna 1
31028 säkerhetsövningar 1
31029 säkerligen 23
31030 säkerställa 55
31031 säkerställande 1
31032 säkerställandet 2
31033 säkerställas 1
31034 säkerställd 1
31035 säkerställer 12
31036 säkerställs 1
31037 säkerställt 1
31038 säkert 62
31039 säkerthetsnormer 1
31040 säkra 43
31041 säkrad 3
31042 säkrade 2
31043 säkrandet 3
31044 säkrar 3
31045 säkrare 4
31046 säkras 3
31047 säkraste 5
31048 säkrat 1
31049 sälja 10
31050 säljare 3
31051 säljas 7
31052 säljer 4
31053 säljförbud 1
31054 säljs 1
31055 säljstart 1
31056 sällan 9
31057 sällsamheter 1
31058 sällsamma 1
31059 sällskap 5
31060 sällskapliga 1
31061 sällskaplighet 1
31062 sällsynt 3
31063 sämre 20
31064 sämst 8
31065 sämsta 1
31066 sända 12
31067 sändas 3
31068 sände 3
31069 sändebud 10
31070 sändebudet 4
31071 sänder 3
31072 sändes 2
31073 sändningar 1
31074 sändningarna 1
31075 sändningsläge 1
31076 sänds 3
31077 säng 3
31078 sängen 7
31079 sängkammare 1
31080 sängkläderna 1
31081 sängs 1
31082 sängöverkastet 1
31083 sänka 14
31084 sänkan 1
31085 sänkas 3
31086 sänker 1
31087 sänkning 3
31088 sänkningar 1
31089 sänkningen 2
31090 sänks 1
31091 sänkt 1
31092 sänkta 1
31093 sänkte 3
31094 sänkts 1
31095 sänt 2
31096 sär 1
31097 särart 1
31098 särarten 1
31099 särarter 1
31100 särbehandla 1
31101 särbehandling 6
31102 särbestämmelse 1
31103 särbestämmelser 1
31104 särdrag 9
31105 särdragen 1
31106 säreget 1
31107 säregna 1
31108 särintressen 2
31109 särkilt 1
31110 särläkemedel 1
31111 särskild 46
31112 särskilda 54
31113 särskilja 2
31114 särskilt 378
31115 säsong 2
31116 säsongsarbete 1
31117 säsongsarbetslöshet 1
31118 säsongsbetonad 1
31119 säsongsbetonade 1
31120 säsongsbundna 2
31121 säsongsjobb 1
31122 säte 4
31123 säten 1
31124 sätet 2
31125 sätt 701
31126 sätta 93
31127 sättandes 1
31128 sättas 14
31129 sätten 3
31130 sätter 36
31131 sättet 71
31132 sätts 14
31133 sättstycken 1
31134 sävliga 1
31135 så 1790
31136 sådan 202
31137 sådana 139
31138 sådant 146
31139 såg 112
31140 såga 1
31141 sågs 2
31142 sågspån 1
31143 sågverk 1
31144 såhär 2
31145 såld 1
31146 sålde 4
31147 såldes 1
31148 således 131
31149 såll 3
31150 sållas 1
31151 sålt 1
31152 sålts 1
31153 sålunda 10
31154 sån 9
31155 såna 7
31156 sång 1
31157 sången 1
31158 sångens 1
31159 sånger 1
31160 sångerna 1
31161 sånt 2
31162 sår 1
31163 såra 1
31164 sårade 2
31165 sårbar 2
31166 sårbara 8
31167 sårbarhet 1
31168 sårbarheten 1
31169 såsom 104
31170 såtillvida 2
31171 såvida 7
31172 såvitt 2
31173 såväl 122
31174 söder 24
31175 söderut 2
31176 södra 26
31177 sögs 1
31178 söka 16
31179 sökande 4
31180 sökanden 1
31181 sökandet 4
31182 sökas 2
31183 söker 25
31184 sökningen 1
31185 sökt 1
31186 sökte 5
31187 sökväg 5
31188 sökvägen 1
31189 sömn 5
31190 söndags 1
31191 söndagstidningar 1
31192 sönder 10
31193 sönderdela 2
31194 sönderdelas 1
31195 sönderdelning 1
31196 sönderdelningsanläggningarna 1
31197 sönderfall 2
31198 söndergrävd 1
31199 sönderklippta 1
31200 sönderrivna 1
31201 sönderslaget 1
31202 sönderslagna 1
31203 sönderslitet 1
31204 söner 4
31205 sörja 10
31206 sörjde 2
31207 sörjer 6
31208 söt 1
31209 söta 1
31210 sötpapper 1
31211 sötvatten 1
31212 sötvattenmatros 1
31213 t 2
31214 t. 1
31215 t.ex 6
31216 t.ex. 59
31217 t.o.m. 18
31218 ta 658
31219 tabell 5
31220 tabellen 3
31221 tabeller 6
31222 tabellerna 2
31223 tabletter 1
31224 tabu 1
31225 tabubelagda 1
31226 tabubelagt 1
31227 tack 92
31228 tacka 178
31229 tackar 58
31230 tacklas 1
31231 tacknämligt 2
31232 tackor 1
31233 tacksam 23
31234 tacksamhet 2
31235 tacksamhetens 1
31236 tacksamma 5
31237 tacksamt 1
31238 tag 20
31239 tagen 3
31240 taget 55
31241 tagg 1
31242 taggar 2
31243 taggarna 2
31244 taggtrådsstaketet 1
31245 tagit 124
31246 tagits 37
31247 tagna 2
31248 tak 8
31249 taken 1
31250 taket 14
31251 takt 14
31252 takten 5
31253 takter 1
31254 taktik 7
31255 taktiska 2
31256 taktiskt 1
31257 taktlöshet 1
31258 takåsarna 1
31259 tal 50
31260 tala 162
31261 talade 82
31262 talades 4
31263 talan 3
31264 talande 2
31265 talang 1
31266 talanger 2
31267 talar 160
31268 talare 37
31269 talaren 11
31270 talares 1
31271 talarlistan 1
31272 talarna 13
31273 talarnas 1
31274 talarstolen 1
31275 talartid 8
31276 talartiden 3
31277 talartiderna 2
31278 talas 29
31279 talat 50
31280 talats 2
31281 talen 2
31282 talesman 5
31283 talesmannen 1
31284 talesmän 1
31285 talesätt 1
31286 talesättet 1
31287 talet 6
31288 talförmågan 1
31289 tallar 1
31290 tallitkatan 1
31291 tallrik 4
31292 tallrikar 1
31293 tallrikarna 1
31294 tallriken 3
31295 tallöst 1
31296 talman 1140
31297 talmannen 11
31298 talmannens 2
31299 talmans 2
31300 talmanskonferens 1
31301 talmanskonferensen 15
31302 talmanskonferensens 1
31303 talmanskonferenser 1
31304 talmän 2
31305 talrika 6
31306 tals 3
31307 tampas 2
31308 tandborste 1
31309 tandem 1
31310 tandlöst 1
31311 tangera 1
31312 tank- 1
31313 tankar 33
31314 tankarna 15
31315 tankbåtar 1
31316 tankbåtarna 2
31317 tanke 151
31318 tankearbetet 1
31319 tankebanor 1
31320 tankefrihet 1
31321 tankegångar 2
31322 tankegångarna 2
31323 tankemöda 1
31324 tanken 40
31325 tankens 1
31326 tankepolis 1
31327 tankern 1
31328 tankerägarnas 1
31329 tankespår 1
31330 tankfartyg 7
31331 tankfartygens 1
31332 tankfartyget 3
31333 tankfordon 1
31334 tankfull 1
31335 tanklöshet 1
31336 tanklöst 1
31337 tankrengöring 2
31338 tankrengöringar 1
31339 tankrengöringarna 1
31340 tant 1
31341 tapeten 2
31342 tappa 6
31343 tappade 2
31344 tappar 3
31345 tappas 1
31346 tappat 2
31347 tappert 1
31348 tappt 1
31349 tar 223
31350 tarifferna 1
31351 tarvligheter 2
31352 tas 132
31353 task 1
31354 tatuerat 1
31355 tavlor 2
31356 tavlorna 1
31357 tax-free 1
31358 tax-free-försäljningen 1
31359 tax-free-lobbyister 1
31360 taxa 1
31361 taxeringsnormer 1
31362 taxi 3
31363 taxichaufför 1
31364 taxifolia 1
31365 taxin 2
31366 taxor 1
31367 taxorna 1
31368 tayloristiska 1
31369 te 7
31370 teater 1
31371 teaterföreställning 1
31372 teatergrupper 1
31373 tecken 27
31374 teckenstorlek 1
31375 tecknade 1
31376 tecknas 1
31377 tecknats 1
31378 tecknen 1
31379 tedde 2
31380 tegel 2
31381 tegeldamm 1
31382 tegelskärva 1
31383 tegelväggen 1
31384 teknik 25
31385 tekniken 16
31386 teknikens 2
31387 tekniker 8
31388 teknikerna 6
31389 teknisk 38
31390 teknisk-ekonomiskt 1
31391 tekniska 88
31392 tekniskt 26
31393 teknokraternas 1
31394 teknologi 3
31395 teknologiska 1
31396 telefon 7
31397 telefonavlyssning 4
31398 telefonavlyssningen 1
31399 telefonbolaget 1
31400 telefonen 2
31401 telefoner 2
31402 telefoni 1
31403 telefonicentren 1
31404 telefonisterna 1
31405 telefonitjänster 1
31406 telefonnummer 1
31407 telefonsamtal 4
31408 telefonsamtalet 2
31409 teleföretagen 1
31410 telegram 2
31411 telekommunikation 4
31412 telekommunikationen 1
31413 telekommunikationer 2
31414 telekommunikationernas 1
31415 telekommunikationsministern 1
31416 telekommunikationsområdet 1
31417 telekommunikationspriserna 1
31418 telekommunikationssektorn 1
31419 telenät 1
31420 teleskop 1
31421 teletrafiken 2
31422 televerket 1
31423 television 1
31424 televisionen 3
31425 televisionsprogrammen 1
31426 tema 1
31427 temat 1
31428 tematisk 2
31429 tematiska 4
31430 tempel 1
31431 temperatur 2
31432 temperaturen 3
31433 temperaturer 4
31434 temperaturhöjningar 1
31435 tempererad 1
31436 tempo 3
31437 temporär 2
31438 temporärt 1
31439 tempot 1
31440 tendens 11
31441 tendensen 9
31442 tendenser 2
31443 tendenserna 3
31444 tendentiöst 1
31445 tenderar 9
31446 tennisbollar 1
31447 tennisskor 1
31448 teokratiskt 1
31449 teologerna 1
31450 teologi 1
31451 teoretisk 2
31452 teoretiska 2
31453 teoretiskt 8
31454 teori 4
31455 teorier 1
31456 teorin 4
31457 ter 1
31458 teratogena 1
31459 teratogent 1
31460 term 2
31461 termen 3
31462 termer 9
31463 termerna 1
31464 terminaler 1
31465 terminen 1
31466 terminis 2
31467 terminologi 1
31468 termins- 1
31469 terminskontrakt 2
31470 territorialitetsprincipen 1
31471 territorialklausul 1
31472 territorialklausulen 3
31473 territorialvatten 1
31474 territorieklausulen 1
31475 territoriell 2
31476 territoriella 15
31477 territorier 5
31478 territoriet 8
31479 territoriets 1
31480 territorium 30
31481 terror 2
31482 terrorbomb 1
31483 terrorism 3
31484 terrorismen 2
31485 terroristattack 2
31486 terroristbomber 1
31487 terrorister 7
31488 terroristerna 2
31489 terroristhandlingar 1
31490 terroristmassaker 1
31491 terrorstyrka 1
31492 terräng 2
31493 terrängen 2
31494 tesen 2
31495 teservis 1
31496 testa 2
31497 testcentrer 1
31498 tester 1
31499 testet 1
31500 teve 1
31501 text 53
31502 text- 1
31503 texten 52
31504 textens 1
31505 texter 11
31506 texterna 5
31507 texternas 1
31508 textilsektorn 1
31509 textredigerare 2
31510 textändring 1
31511 that 1
31512 thatcherianska 1
31513 the 28
31514 therefore 1
31515 tibetaner 1
31516 tibetanerna 3
31517 tibetanska 5
31518 tid 217
31519 tiden 155
31520 tidens 6
31521 tider 14
31522 tiderna 1
31523 tidevarv 2
31524 tidig 5
31525 tidiga 9
31526 tidigare 228
31527 tidigarelagda 1
31528 tidigareläggas 1
31529 tidigt 26
31530 tidlöshet 1
31531 tidning 3
31532 tidningar 5
31533 tidningarna 2
31534 tidningen 7
31535 tidningsartikel 2
31536 tidningsintervju 1
31537 tidningsreferat 1
31538 tidplanen 1
31539 tidpunkt 22
31540 tidpunkten 10
31541 tidpunkter 1
31542 tids 4
31543 tidsaspekt 1
31544 tidsbegränsade 1
31545 tidsbegränsningen 3
31546 tidsbestämda 2
31547 tidsbestämmas 1
31548 tidsbrist 2
31549 tidsfaktorn 1
31550 tidsfrist 10
31551 tidsfristen 6
31552 tidsfristens 1
31553 tidsfrister 9
31554 tidsfält 1
31555 tidsglappet 1
31556 tidsgräns 1
31557 tidshorisont 1
31558 tidsinställd 2
31559 tidskontrakt 1
31560 tidsmässiga 2
31561 tidsperiod 6
31562 tidsperioder 1
31563 tidsplan 9
31564 tidsplanen 7
31565 tidspress 1
31566 tidsproblematiken 1
31567 tidsram 1
31568 tidsramar 5
31569 tidsramarna 2
31570 tidsramen 1
31571 tidsrymd 3
31572 tidsrymden 1
31573 tidsschemat 2
31574 tidsskede 1
31575 tidsskäl 1
31576 tidsskänken 1
31577 tidsålder 2
31578 tidsåtgång 1
31579 tidsödande 1
31580 tidtabell 17
31581 tidtabellen 2
31582 tidvatten 3
31583 tidvattnet 1
31584 tiga 2
31585 tigande 1
31586 tiger 5
31587 tigern 1
31588 tiggde 1
31589 tigger 1
31590 till 6113
31591 tillade 5
31592 tillagades 1
31593 tillbad 1
31594 tillbaka 189
31595 tillbakablick 1
31596 tillbakadragande 2
31597 tillbakadragandet 2
31598 tillbakadragen 1
31599 tillbakadragna 1
31600 tillbakagång 13
31601 tillbakalutad 1
31602 tillbakavisa 3
31603 tillbakavisande 2
31604 tillbakavisar 5
31605 tillbakavisat 1
31606 tillbakavisats 2
31607 tillbaks 4
31608 tillbehör 1
31609 tillblivelse 1
31610 tillbringa 3
31611 tillbringade 1
31612 tillbringat 3
31613 tillbud 1
31614 tillbörligt 1
31615 tilldela 2
31616 tilldelad 1
31617 tilldelade 1
31618 tilldelades 4
31619 tilldelar 2
31620 tilldelas 7
31621 tilldelats 7
31622 tilldelning 5
31623 tilldelningen 2
31624 tilldragelse 1
31625 tillerkände 1
31626 tillerkänner 3
31627 tillerkänns 1
31628 tillfalla 1
31629 tillfaller 1
31630 tillfinnandes 1
31631 tillflyktsort 1
31632 tillfoga 7
31633 tillfogar 1
31634 tillfogat 1
31635 tillfogats 1
31636 tillfreds 3
31637 tillfredsställa 4
31638 tillfredsställande 29
31639 tillfredsställde 1
31640 tillfredsställelse 14
31641 tillfrågad 1
31642 tillfrågats 1
31643 tillfälle 69
31644 tillfällen 41
31645 tillfället 32
31646 tillfällig 7
31647 tillfälliga 8
31648 tillfällighet 11
31649 tillfälligheter 1
31650 tillfälligt 12
31651 tillfälligtvis 1
31652 tillfångatagande 1
31653 tillför 9
31654 tillföra 8
31655 tillföras 1
31656 tillförlitlig 3
31657 tillförlitliga 4
31658 tillförlitlighet 2
31659 tillförlitlighetsproblem 1
31660 tillförlitligt 2
31661 tillförordnad 2
31662 tillförs 1
31663 tillförsikt 5
31664 tillförsäkra 1
31665 tillförsäkrar 1
31666 tillfört 1
31667 tillgivenhet 4
31668 tillgivet 1
31669 tillgodoräkna 1
31670 tillgodose 4
31671 tillgodosedda 2
31672 tillgodoser 1
31673 tillgodoses 3
31674 tillgripa 3
31675 tillgripas 1
31676 tillgriper 2
31677 tillgänglig 15
31678 tillgängliga 47
31679 tillgänglighet 3
31680 tillgängligheten 3
31681 tillgängligt 8
31682 tillgå 2
31683 tillgång 78
31684 tillgångar 10
31685 tillgången 18
31686 tillhandahålla 33
31687 tillhandahållande 25
31688 tillhandahållandet 2
31689 tillhandahållas 5
31690 tillhandahåller 12
31691 tillhandahållit 2
31692 tillhandahållits 5
31693 tillhandahållna 1
31694 tillhandahålls 3
31695 tillhandahöll 2
31696 tillhåll 1
31697 tillhör 31
31698 tillhöra 6
31699 tillhörande 2
31700 tillhörde 5
31701 tillhörighet 2
31702 tillhörigheten 2
31703 tillhörigheter 2
31704 tillika 3
31705 tillintetgjorts 1
31706 tillintetgöra 1
31707 tillit 2
31708 tillkom 3
31709 tillkommande 1
31710 tillkommer 9
31711 tillkommit 5
31712 tillkomst 2
31713 tillkomsten 1
31714 tillkrånglade 1
31715 tillkännagav 4
31716 tillkännage 2
31717 tillkännager 7
31718 tillkännages 3
31719 tillkännagett 1
31720 tillkännagivanden 3
31721 tillkännagivandena 1
31722 tillkännagivit 2
31723 tillkännagivits 1
31724 tillkännagivna 1
31725 tillmätas 1
31726 tillmäter 2
31727 tillmäts 2
31728 tillmötes 1
31729 tillmötesgå 2
31730 tillmötesgående 4
31731 tillmötesgås 1
31732 tillmötesgått 1
31733 tillnärmelsevis 1
31734 tillnärmning 11
31735 tillnärmningen 1
31736 tillnärmningsprocess 1
31737 tillrop 1
31738 tillryggalagt 1
31739 tillryggalagts 1
31740 tillryggalägger 1
31741 tillräcklig 39
31742 tillräckliga 17
31743 tillräckligt 115
31744 tillrätta 2
31745 tillrättalägger 1
31746 tillrättavisare 1
31747 tillrådligt 1
31748 tills 34
31749 tillsammans 152
31750 tillsats 3
31751 tillsatsdirektivet 1
31752 tillsatser 18
31753 tillsatserna 3
31754 tillsatsernas 1
31755 tillsatsämnen 1
31756 tillsatt 2
31757 tillsattes 1
31758 tillsatts 1
31759 tillse 13
31760 tillskansa 2
31761 tillskansar 1
31762 tillskapade 1
31763 tillskapandet 1
31764 tillskott 6
31765 tillskriver 2
31766 tillskrivs 1
31767 tillskyndar 2
31768 tillsluta 1
31769 tillstymmelse 1
31770 tillställa 1
31771 tillställningar 1
31772 tillställningarna 2
31773 tillställningen 2
31774 tillstå 2
31775 tillstånd 35
31776 tillstånden 2
31777 tillståndet 9
31778 tillståndsförfarandena 1
31779 tillståndssystem 1
31780 tillstår 1
31781 tillstås 1
31782 tillsyn 4
31783 tillsynsmyndighetens 1
31784 tillsynsmyndigheter 1
31785 tillsätt 1
31786 tillsätta 3
31787 tillsättandet 2
31788 tillsätter 1
31789 tillsättning 1
31790 tillsättningar 1
31791 tillsätts 3
31792 tillta 1
31793 tilltagande 2
31794 tilltal 1
31795 tilltala 1
31796 tilltalade 2
31797 tilltalande 1
31798 tilltalar 3
31799 tilltar 1
31800 tilltro 2
31801 tilltron 1
31802 tillträdandet 1
31803 tillträdde 1
31804 tillträde 29
31805 tillträdet 4
31806 tilltänkta 1
31807 tillval 1
31808 tillvara 3
31809 tillvarata 1
31810 tillvaro 8
31811 tillvaron 2
31812 tillverka 5
31813 tillverkade 2
31814 tillverkar 3
31815 tillverkaransvar 1
31816 tillverkaransvaret 4
31817 tillverkare 3
31818 tillverkaren 11
31819 tillverkarens 2
31820 tillverkarna 15
31821 tillverkarnas 6
31822 tillverkas 4
31823 tillverkats 2
31824 tillverkning 3
31825 tillverkningen 4
31826 tillverkningsindustri 1
31827 tillverkningsindustrin 5
31828 tillverkningsprocesser 1
31829 tillverkningssektorn 2
31830 tillväga 6
31831 tillvägagångssätt 23
31832 tillvägagångssätten 1
31833 tillvägagångssättet 4
31834 tillväxt 78
31835 tillväxt- 2
31836 tillväxtbefrämjande 1
31837 tillväxtbranscherna 1
31838 tillväxtcentrum 1
31839 tillväxtdynamik 1
31840 tillväxten 30
31841 tillväxtfaktor 1
31842 tillväxtfaktorer 1
31843 tillväxtmål 2
31844 tillväxtmålsättningar 1
31845 tillväxtnivå 4
31846 tillväxtnivåer 1
31847 tillväxtpotential 1
31848 tillväxtprognosen 1
31849 tillväxttakt 2
31850 tillväxtökande 1
31851 tillägg 15
31852 tillägga 21
31853 tillägget 1
31854 tilläggs 1
31855 tilläggsbudget 1
31856 tilläggsfråga 3
31857 tilläggskrav 1
31858 tillägna 2
31859 tillämpa 83
31860 tillämpad 1
31861 tillämpade 1
31862 tillämpades 1
31863 tillämpande 1
31864 tillämpandet 1
31865 tillämpar 16
31866 tillämpas 93
31867 tillämpat 2
31868 tillämpats 9
31869 tillämplig 7
31870 tillämpliga 9
31871 tillämplighet 2
31872 tillämpligt 4
31873 tillämpning 63
31874 tillämpningar 1
31875 tillämpningarna 1
31876 tillämpningen 61
31877 tillämpningsbestämmelser 1
31878 tillämpningsbestämmelserna 2
31879 tillämpningsförfaranden 1
31880 tillämpningsförordning 1
31881 tillämpningsförordningen 2
31882 tillämpningsområde 6
31883 tillämpningsområdet 6
31884 tillämpningsprocessen 1
31885 tillämpningsstrategier 1
31886 tillämpningssvårigheter 1
31887 tillämpningsövervakning 1
31888 tillät 1
31889 tillåt 2
31890 tillåta 35
31891 tillåtande 1
31892 tillåtas 13
31893 tillåtelse 1
31894 tillåten 6
31895 tillåter 50
31896 tillåtet 5
31897 tillåtits 1
31898 tillåtliga 1
31899 tillåtna 12
31900 tillåts 11
31901 timing 1
31902 timjan 1
31903 timma 1
31904 timmar 28
31905 timmarna 1
31906 timmars 1
31907 timme 15
31908 ting 21
31909 tingens 1
31910 tinninglockar 2
31911 tinningådror 1
31912 tio 56
31913 tionde 1
31914 tionyheterna 1
31915 tiopundssedlarna 1
31916 tiotal 3
31917 tiotals 8
31918 tiotusen 1
31919 tiotusentals 5
31920 tioåriga 1
31921 tioårsperioden 1
31922 tips 2
31923 tipsade 1
31924 tisdag 3
31925 tisdagen 3
31926 tisdagens 1
31927 titan 1
31928 titel 2
31929 titeln 11
31930 titelsektionen 1
31931 titelsidan 1
31932 titlar 1
31933 titt 7
31934 titta 57
31935 tittade 34
31936 tittande 2
31937 tittar 20
31938 tittarnöje 1
31939 tja 1
31940 tjata 1
31941 tjatig 1
31942 tjeckiske 2
31943 tjejer 1
31944 tjetjenska 4
31945 tjetjenskt 2
31946 tjock 4
31947 tjocka 6
31948 tjockisen 1
31949 tjockleken 1
31950 tjockolja 2
31951 tjugo 11
31952 tjugofem 5
31953 tjugoförsta 2
31954 tjugonde 4
31955 tjugosex 2
31956 tjugosexåriga 1
31957 tjugosju 2
31958 tjugotusen 2
31959 tjugotvå 1
31960 tjugotvåtusen 1
31961 tjugu 1
31962 tjur 1
31963 tjuren 2
31964 tjurskallig 1
31965 tjusade 1
31966 tjusar 1
31967 tjusat 1
31968 tjusig 2
31969 tjusning 1
31970 tjuvnad 1
31971 tjäna 14
31972 tjänade 1
31973 tjänar 26
31974 tjänare 2
31975 tjänaren 1
31976 tjänarstaben 1
31977 tjänas 1
31978 tjänat 6
31979 tjänst 35
31980 tjänstberett 1
31981 tjänsteenhet 1
31982 tjänsteenheter 4
31983 tjänsteenheterna 1
31984 tjänstefel 1
31985 tjänsteföreskrifterna 6
31986 tjänsteföretag 1
31987 tjänsteföretagen 2
31988 tjänstekriterier 1
31989 tjänstekvaliteten 3
31990 tjänsteleverantören 2
31991 tjänsteman 9
31992 tjänstemanna-apparaten 1
31993 tjänstemannakårer 1
31994 tjänstemannarepresentanter 1
31995 tjänstemän 42
31996 tjänstemännen 11
31997 tjänstemännens 4
31998 tjänstemäns 3
31999 tjänsten 6
32000 tjänstenivå 5
32001 tjänstenivån 2
32002 tjänstens 1
32003 tjänsteproducenter 3
32004 tjänsteproducenterna 1
32005 tjänsteproducenters 1
32006 tjänsteproduktion 1
32007 tjänster 111
32008 tjänsterna 22
32009 tjänsternas 1
32010 tjänsterum 1
32011 tjänstesektorer 1
32012 tjänstesektorn 4
32013 tjänsteuppdrag 2
32014 tjänsteutbudet 1
32015 tjänsteåligganden 1
32016 tjänstgjorde 1
32017 tjänstgjort 1
32018 tjänstgör 1
32019 tjänstgörande 15
32020 tjära 2
32021 tjöt 1
32022 to 2
32023 toalettbord 1
32024 toaletten 3
32025 toaletter 1
32026 toaletterna 2
32027 toalettköerna 1
32028 tobak 2
32029 tobaksblommorna 1
32030 tobaksodling 1
32031 tobakspung 1
32032 toddyn 1
32033 todo 1
32034 tofflor 2
32035 tofflorna 1
32036 tofsar 1
32037 tog 128
32038 toga 1
32039 togorna 1
32040 togs 25
32041 tokig 2
32042 tolerans 15
32043 toleransen 1
32044 toleranskulturen 1
32045 tolerant 1
32046 toleranta 3
32047 tolerera 3
32048 tolererar 1
32049 tolereras 7
32050 tolk 1
32051 tolka 8
32052 tolkade 3
32053 tolkar 10
32054 tolkarna 4
32055 tolkarnas 1
32056 tolkas 13
32057 tolkat 1
32058 tolkats 2
32059 tolkning 20
32060 tolkningar 4
32061 tolkningarna 1
32062 tolkningarnas 1
32063 tolkningen 11
32064 tolkningsmeddelanden 1
32065 tolkningsmöjligheterna 1
32066 tolkningsproblem 1
32067 tolv 9
32068 tom 6
32069 tomater 3
32070 tomatkonserver 1
32071 tomatpuré 1
32072 tomhet 3
32073 tomma 11
32074 tomrum 5
32075 tomtarna 1
32076 ton 35
32077 toner 1
32078 tonfall 4
32079 tonfisk 18
32080 tonfiskbestånden 1
32081 tonfisken 5
32082 tonfisket 1
32083 tonfiskliknande 1
32084 tongivande 1
32085 tongångar 1
32086 tonlös 1
32087 tonvikt 6
32088 tonvikten 3
32089 tonåringar 2
32090 tonårsgrammofonen 1
32091 topp 4
32092 toppen 8
32093 toppluva 1
32094 toppmöte 14
32095 toppmöten 3
32096 toppmötena 1
32097 toppmötesnivå 1
32098 toppmötet 73
32099 toppnyhet 1
32100 toppositioner 1
32101 topprioritet 1
32102 topptjänstemän 1
32103 torde 5
32104 tordönsröst 1
32105 torftig 1
32106 torg 1
32107 torka 12
32108 torkade 3
32109 torkan 1
32110 torkas 1
32111 torkat 1
32112 torna 1
32113 tornet 1
32114 torniga 1
32115 torpet 2
32116 torra 4
32117 torrare 1
32118 torrhet 1
32119 torrlägger 1
32120 torrt 2
32121 torsdag 15
32122 torsdagen 7
32123 torsdagens 1
32124 torsdags 1
32125 torsk 3
32126 torskbestånden 1
32127 torsken 1
32128 torskfiske 1
32129 torskkvot 1
32130 torskkvoten 1
32131 torteras 2
32132 torterats 1
32133 tortyr 4
32134 tortyren 1
32135 tortyrinstrument 1
32136 torven 4
32137 torvvatten 1
32138 total 14
32139 totala 35
32140 totalanslag 2
32141 totalanslaget 3
32142 totalansvar 1
32143 totalbeloppet 1
32144 totalblockad 1
32145 totalfångst 2
32146 totalfångsten 2
32147 totalförbud 2
32148 totalförstört 1
32149 totalitarism 2
32150 totalitarismens 1
32151 totalitära 2
32152 totalsumma 1
32153 totalsumman 1
32154 totalt 22
32155 totalvolym 1
32156 toxiska 1
32157 trader 1
32158 tradition 15
32159 traditionalism 1
32160 traditionell 4
32161 traditionella 16
32162 traditionellt 4
32163 traditionen 6
32164 traditionens 1
32165 traditioner 8
32166 traditionerna 2
32167 trafik 5
32168 trafik- 1
32169 trafikanter 1
32170 trafikeländet 1
32171 trafiken 7
32172 trafikens 1
32173 trafikerar 1
32174 trafikkontroller 1
32175 trafikled 1
32176 trafikolyckor 1
32177 trafikpolisen 1
32178 trafikpoliser 1
32179 trafikstockningar 1
32180 trafiksäkerhet 1
32181 trafiksäkerheten 8
32182 trafikön 1
32183 tragedi 10
32184 tragedier 6
32185 tragedin 6
32186 tragisk 4
32187 tragiska 12
32188 tragiskt 8
32189 trakasserad 1
32190 trakasserier 3
32191 trakt 1
32192 trakten 1
32193 trakterna 1
32194 tramp 2
32195 trampar 1
32196 trans 3
32197 transaktioner 2
32198 transaktionskostnader 1
32199 transatlantiska 2
32200 transeuropeiska 7
32201 transferable 2
32202 transfereringar 1
32203 transformera 2
32204 transformeras 3
32205 transithallen 1
32206 transitivt 1
32207 transitland 2
32208 transitländer 1
32209 transitrutten 1
32210 transittrafiken 1
32211 transmissibel 1
32212 transnationell 3
32213 transnationella 6
32214 transnationellt 4
32215 transparens 1
32216 transparent 1
32217 transport 78
32218 transport- 5
32219 transportabla 1
32220 transportbeställarna 1
32221 transportbestämmelser 1
32222 transportdirektiv 1
32223 transporten 7
32224 transporter 27
32225 transportera 3
32226 transporterade 2
32227 transporterades 1
32228 transporterar 2
32229 transporteras 8
32230 transporterna 5
32231 transportfederationen 1
32232 transportfrågor 1
32233 transportgruppen 1
32234 transportkapacitet 1
32235 transportkostnaderna 2
32236 transportmarknad 1
32237 transportmedel 1
32238 transportministrar 1
32239 transportnät 3
32240 transportnäten 2
32241 transportområden 1
32242 transportområdet 2
32243 transportpolitik 1
32244 transportpolitiken 2
32245 transportpolitiker 1
32246 transportpolitiska 1
32247 transportproblem 1
32248 transportsektorn 2
32249 transportsäkerhet 3
32250 transportsäkerheten 3
32251 transportsätt 1
32252 transportutskottet 1
32253 transportörernas 1
32254 trappa 2
32255 trappan 11
32256 trappavsatsen 2
32257 trapphallen 1
32258 trapporna 1
32259 trappsteg 1
32260 trappsteget 1
32261 trasa 1
32262 trasas 1
32263 trasig 3
32264 trasiga 5
32265 trasigt 2
32266 trasmatta 1
32267 trasmattan 1
32268 trasor 1
32269 trassel 1
32270 trassla 1
32271 trasslade 2
32272 trasslat 1
32273 trasslig 1
32274 tratt 1
32275 traumatiska 1
32276 travar 3
32277 traven 2
32278 travesterade 1
32279 tre 179
32280 tre-fyra 1
32281 trea 1
32282 trebent 1
32283 tredagarskryssning 1
32284 tredelade 1
32285 tredje 191
32286 tredjedel 12
32287 tredjedelar 4
32288 tredjelandsmedborgare 7
32289 tredjelandsmedborgares 1
32290 trehjulingar 1
32291 trehundrafemti 1
32292 trekilometerspromenad 1
32293 treklang 1
32294 tremånadersfristen 1
32295 tremånadersperioden 2
32296 trend 4
32297 trenden 3
32298 trender 1
32299 trepartsagerande 1
32300 trepartsarbete 1
32301 trepartsarbetsgrupp 3
32302 trepartsarbetsgruppen 1
32303 trepartsmöte 1
32304 trepartssamtalen 1
32305 trephena-mat 1
32306 treprocentsnormen 1
32307 trettio 12
32308 trettiofem 3
32309 trettiofemårsåldern 1
32310 trettiotal 1
32311 trettiotalet 3
32312 trettioåtta 1
32313 tretton 7
32314 trettonde 1
32315 trettonåriga 1
32316 trevlig 3
32317 trevliga 1
32318 trevligt 5
32319 treårsperioder 1
32320 triangel 1
32321 triangelformad 1
32322 triangelförhållande 1
32323 tribunal 2
32324 tribunen 1
32325 tributyl 1
32326 trick 1
32327 trickle 1
32328 trikåfabrik 1
32329 trilby 1
32330 trilbyhatt 1
32331 triljoner 1
32332 trimmade 1
32333 trio 1
32334 trirem 1
32335 trissa 1
32336 trist 5
32337 trista 1
32338 triumf 1
32339 triumferande 1
32340 triumferat 1
32341 trivas 1
32342 trivdes 3
32343 trivialaste 1
32344 trivsamma 1
32345 tro 64
32346 trodde 28
32347 troddes 1
32348 trofasthet 1
32349 troféer 1
32350 trogen 5
32351 troget 2
32352 trogne 1
32353 trojanska 1
32354 trojkan 1
32355 troliga 1
32356 troligen 10
32357 troligt 6
32358 troligtvis 4
32359 trolla 2
32360 trolldom 2
32361 trolldomsböcker 1
32362 trolldomskraft 1
32363 trolleri 1
32364 trolleriet 1
32365 trollformler 1
32366 trollguld 1
32367 trollkarl 5
32368 trollkarlar 5
32369 trollkarlen 1
32370 trollkarlsbutik 1
32371 trollkarlshatt 1
32372 trollkarlshem 1
32373 trollkarlsskolan 1
32374 trollkarlsvärlden 4
32375 trollkonst 1
32376 trollspö 3
32377 trollspöt 1
32378 trollstav 3
32379 trollstaven 1
32380 tron 1
32381 tropikerna 1
32382 tropisk 1
32383 tropiska 15
32384 tror 487
32385 trosartikel 1
32386 trots 155
32387 trott 7
32388 trottoaren 2
32389 trottoarer 1
32390 trottoarerna 1
32391 trovärdig 8
32392 trovärdiga 8
32393 trovärdige 1
32394 trovärdighet 29
32395 trovärdigheten 4
32396 trovärdighetskris 1
32397 trovärdighetsproblem 1
32398 trovärdighetstest 1
32399 trovärdighetstestet 1
32400 trovärdigt 2
32401 trubbigt 1
32402 trumfkort 3
32403 trummade 1
32404 trummorna 1
32405 trumpet 1
32406 trumpinnar 1
32407 trupper 8
32408 truppminor 1
32409 trusten 1
32410 truster 2
32411 trusterna 1
32412 tryck 15
32413 trycka 7
32414 tryckalster 1
32415 tryckas 2
32416 tryckbärande 1
32417 trycker 2
32418 trycket 8
32419 tryckfel 1
32420 tryckfriheten 1
32421 tryckningen 1
32422 tryckta 2
32423 tryckte 6
32424 trygg 1
32425 trygga 3
32426 tryggad 1
32427 tryggande 1
32428 tryggas 1
32429 trygghet 52
32430 tryggheten 37
32431 trygghetsmodellen 1
32432 trygghetsnivå 1
32433 trygghetspolitik 1
32434 trygghetssystem 9
32435 trygghetssystemen 21
32436 trygghetssystemens 3
32437 trygghetssystemet 4
32438 tryggt 3
32439 trä 4
32440 träbord 1
32441 träd 12
32442 träda 19
32443 trädde 13
32444 träddungar 1
32445 träddunge 1
32446 träden 9
32447 träder 12
32448 trädet 1
32449 trädgård 2
32450 trädgårdar 2
32451 trädgården 8
32452 trädgårdsanläggningarna 1
32453 trädgårdsbänken 3
32454 trädgårdshäcken 1
32455 trädgårdsmöbeln 1
32456 trädgårdsprodukter 1
32457 trädgårdsstolarna 1
32458 trädstruktur 1
32459 trädtopparna 1
32460 träffa 16
32461 träffade 14
32462 träffades 4
32463 träffande 3
32464 träffar 7
32465 träffas 10
32466 träffat 2
32467 träffats 3
32468 träkolsgrill 1
32469 träldom 2
32470 trälåda 1
32471 tränat 1
32472 tränga 2
32473 trängande 1
32474 trängda 1
32475 trängde 6
32476 trängdes 1
32477 tränger 4
32478 trängt 2
32479 träning 1
32480 träproduktion 1
32481 träsk 2
32482 träskulpturerna 1
32483 träskylt 1
32484 trätor 1
32485 trätt 10
32486 tråd 4
32487 trådar 4
32488 trådarna 1
32489 trådbar 1
32490 trådde 1
32491 tråden 2
32492 tråkigaste 1
32493 tråkigt 8
32494 trålar 1
32495 trånga 1
32496 trångmål 1
32497 trångt 2
32498 tröga 2
32499 tröghet 5
32500 trögheten 2
32501 tröja 1
32502 tröskade 1
32503 tröskar 1
32504 tröskel 3
32505 tröskeln 5
32506 tröskelvärdet 1
32507 tröst 3
32508 tröstad 1
32509 tröstade 1
32510 tröstegrund 1
32511 trött 6
32512 trötta 3
32513 trötthet 3
32514 tröttheten 1
32515 tröttnade 2
32516 tröttsamma 1
32517 tröttsamt 1
32518 tsetseflugor 1
32519 tudelad 1
32520 tuff 1
32521 tuffare 1
32522 tuffingarna 1
32523 tufft 2
32524 tuggummi 1
32525 tuggummit 1
32526 tull 2
32527 tull- 1
32528 tullavgifter 1
32529 tullavgifterna 1
32530 tullförvaltningen 1
32531 tullgåvor 1
32532 tullhinder 1
32533 tullhus 1
32534 tullintegration 1
32535 tullkontroll 1
32536 tullmyndighet 1
32537 tullmyndigheten 1
32538 tullmyndigheter 1
32539 tullmyndigheterna 3
32540 tullsamarbetskommittén 1
32541 tulltariff 1
32542 tulltjänstemän 2
32543 tulltjänstemännen 1
32544 tulltjänstemännens 1
32545 tulltjänster 1
32546 tullättnader 1
32547 tum 1
32548 tumma 3
32549 tummarna 1
32550 tummen 1
32551 tumultet 1
32552 tumultuarisk 1
32553 tunc 1
32554 tung 15
32555 tunga 13
32556 tungmetaller 8
32557 tungmetallerna 1
32558 tungrodd 1
32559 tungrodda 1
32560 tungroddhet 1
32561 tungsint 1
32562 tungt 8
32563 tunn 2
32564 tunna 6
32565 tunnades 1
32566 tunneln 2
32567 tunneltrafik 1
32568 tunnland 2
32569 tunnlar 3
32570 tunnlarna 1
32571 tunt 3
32572 tur 30
32573 turer 1
32574 turism 70
32575 turismen 50
32576 turismens 4
32577 turismfrågor 1
32578 turista 1
32579 turistbranschen 2
32580 turistbyråerna 1
32581 turistcentrer 2
32582 turister 4
32583 turisterna 2
32584 turisthandel 1
32585 turistindustri 1
32586 turistindustrin 6
32587 turistiskt 2
32588 turistland 1
32589 turistmarknaden 3
32590 turistmål 1
32591 turistmålet 1
32592 turistnäring 4
32593 turistnäringen 18
32594 turistnäringens 4
32595 turistområde 1
32596 turistområdet 1
32597 turistorterna 1
32598 turistpolitik 3
32599 turistpolitiken 2
32600 turistpotential 1
32601 turistsektorers 1
32602 turistsektorn 5
32603 turistsäsongen 2
32604 turistutbildningen 1
32605 turkar 2
32606 turkarna 2
32607 turkarnas 1
32608 turkcyprioter 1
32609 turkcyprioterna 1
32610 turkcypriotiska 6
32611 turkcypriotiske 1
32612 turkisk-grekiska 1
32613 turkiska 20
32614 turkiske 3
32615 turkiskt 1
32616 turn-over 1
32617 tusan 2
32618 tusen 17
32619 tusentals 24
32620 tuta 1
32621 tutade 2
32622 tv-sända 1
32623 tv-teknik 1
32624 tveka 5
32625 tvekade 1
32626 tvekan 43
32627 tvekar 8
32628 tvekat 2
32629 tveklöst 4
32630 tveksam 5
32631 tveksamhet 2
32632 tveksamma 2
32633 tveksamt 3
32634 tvetydig 3
32635 tvetydiga 3
32636 tvetydighet 5
32637 tvetydigheten 1
32638 tvetydigheter 1
32639 tvillingarna 1
32640 tvillingbröder 1
32641 tvillingpar 1
32642 tvillingpropeller 1
32643 tvinga 17
32644 tvingad 2
32645 tvingade 6
32646 tvingades 5
32647 tvingande 11
32648 tvingar 15
32649 tvingas 28
32650 tvingats 4
32651 tvinnade 2
32652 tvist 4
32653 tvista 1
32654 tvistefrågor 1
32655 tvisten 1
32656 tvister 6
32657 tvivel 68
32658 tvivelaktig 3
32659 tvivelaktiga 2
32660 tvivelsmålen 1
32661 tvivelsutan 3
32662 tvivla 1
32663 tvivlar 17
32664 tvivlat 1
32665 tvungen 31
32666 tvungna 23
32667 tvärgående 2
32668 tvärpolitiska 2
32669 tvärs 7
32670 tvärsöver 1
32671 tvärt 2
32672 tvärtemot 4
32673 tvärtom 36
32674 tvätta 4
32675 tvättade 2
32676 tvättat 1
32677 tvätten 1
32678 tvättfat 1
32679 tvättmedelseksem 1
32680 två 428
32681 två-ett 1
32682 två-penny-halv-penny 1
32683 två-tre 1
32684 tvåhundra 5
32685 tvåhundraåriga 1
32686 tvålbit 1
32687 tvålen 1
32688 tvålflingor 1
32689 tvång 5
32690 tvånget 3
32691 tvångsarbetarna 2
32692 tvångsfinansieras 1
32693 tvångsförflyttade 2
32694 tvångsförflyttats 2
32695 tvångsintegrerats 1
32696 tvångsmarschen 1
32697 tvångsmedel 1
32698 tvångsmekanism 1
32699 tvångsrekryteras 1
32700 tvångsstruktur 1
32701 tvångströja 1
32702 tvångströjor 1
32703 tvåprocentströskeln 1
32704 tvåspråksutbildningen 1
32705 tvåtusen 1
32706 tvåårig 1
32707 tvååriga 1
32708 twist 1
32709 ty 31
32710 tycka 8
32711 tyckas 3
32712 tycke 4
32713 tycker 197
32714 tycks 33
32715 tyckt 5
32716 tyckte 28
32717 tycktes 19
32718 tyckts 1
32719 tydde 1
32720 tyder 13
32721 tydlig 45
32722 tydliga 44
32723 tydligare 19
32724 tydligaste 3
32725 tydligen 17
32726 tydliggjorde 1
32727 tydliggjort 2
32728 tydliggör 4
32729 tydliggöra 4
32730 tydliggöras 1
32731 tydliggörs 1
32732 tydlighet 10
32733 tydligt 170
32734 tyg 2
32735 tygellösa 1
32736 tygla 1
32737 tygleksaker 1
32738 tynande 1
32739 tynga 2
32740 tyngande 1
32741 tyngas 1
32742 tyngd 7
32743 tyngdpunkt 1
32744 tyngdpunkten 3
32745 tyngdpunkter 1
32746 tynger 3
32747 tyngre 1
32748 tyngst 1
32749 tyngsta 1
32750 typ 77
32751 typen 36
32752 typer 21
32753 typerna 2
32754 typexempel 1
32755 typfall 1
32756 typgodkännanden 1
32757 typisk 1
32758 typiska 1
32759 typiskt 2
32760 typsnitt 1
32761 typtrogen 1
32762 tyranners 1
32763 tyranni 4
32764 tysk 2
32765 tyska 34
32766 tyskar 1
32767 tyskarna 1
32768 tyske 3
32769 tyskspråkig 1
32770 tyskt 2
32771 tyst 19
32772 tysta 7
32773 tystar 1
32774 tystare 2
32775 tystlåten 1
32776 tystlåtne 1
32777 tystnad 14
32778 tystnade 3
32779 tystnaden 2
32780 tystnar 1
32781 tyvärr 79
32782 täcka 6
32783 täckande 1
32784 täckas 2
32785 täcker 18
32786 täckmantel 1
32787 täcks 8
32788 täckt 3
32789 täckte 2
32790 tält 2
32791 tältet 2
32792 tämligen 7
32793 tända 1
32794 tändanordningarna 1
32795 tändas 1
32796 tände 3
32797 tänder 6
32798 tänderna 1
32799 tändes 2
32800 tänds 1
32801 tändsticka 1
32802 tändstickor 2
32803 tänja 1
32804 tänjas 1
32805 tänk 7
32806 tänka 93
32807 tänkande 1
32808 tänkandet 2
32809 tänkas 8
32810 tänkbar 1
32811 tänkbara 9
32812 tänkbart 2
32813 tänker 115
32814 tänkesättet 1
32815 tänkt 15
32816 tänkta 2
32817 tänkte 34
32818 tänktes 1
32819 tänkvärt 1
32820 tänt 1
32821 täppa 4
32822 täpper 1
32823 tärningsspel 1
32824 tärt 2
32825 täta 3
32826 tätare 2
32827 tätbefolkat 2
32828 täten 3
32829 tätortsområden 1
32830 tätt 3
32831 tävla 1
32832 tävlade 1
32833 tävlar 3
32834 tävling 2
32835 tå 5
32836 tåg 5
32837 tåg- 1
32838 tåget 3
32839 tågets 1
32840 tågkraschen 1
32841 tågolyckan 1
32842 tål 1
32843 tålamod 4
32844 tålig 1
32845 tåligt 1
32846 tålmodigt 1
32847 tån 1
32848 tårstrimmiga 1
32849 tårta 2
32850 töckniga 1
32851 töcknigt 1
32852 tömd 1
32853 tömde 1
32854 tömma 1
32855 tömmer 1
32856 töms 4
32857 tömt 1
32858 törnbusken 1
32859 törs 1
32860 u-länderna 4
32861 u-ländernas 1
32862 udda 3
32863 uggla 3
32864 ugglan 2
32865 ugglor 1
32866 ugn 1
32867 ugnen 1
32868 ull 2
32869 ulliga 1
32870 ultimatum 1
32871 ultraliberala 4
32872 ultraliberalism 1
32873 ultraperifer 1
32874 ultraperifera 2
32875 umbärande 1
32876 umgänge 1
32877 umgängesformer 1
32878 umgänget 1
32879 umgås 1
32880 umgåtts 1
32881 un 2
32882 una 2
32883 und 1
32884 undan 28
32885 undanber 2
32886 undandrar 1
32887 undandras 1
32888 undanflykter 2
32889 undanforslad 1
32890 undanglidande 1
32891 undanhålla 2
32892 undanmanövrar 1
32893 undanröja 12
32894 undanröjas 1
32895 undanröjer 1
32896 undanröjts 1
32897 undanslagna 1
32898 undanta 6
32899 undantag 60
32900 undantagen 6
32901 undantaget 6
32902 undantagna 3
32903 undantagsbestämmelser 1
32904 undantagsfall 2
32905 undantagsförfarandet 1
32906 undantagsförordning 1
32907 undantagsmässig 1
32908 undantagsperiod 1
32909 undantagsregeln 3
32910 undantagsregler 1
32911 undantagssituationer 1
32912 undantagstillstånd 1
32913 undantagstillståndet 1
32914 undantagsvis 1
32915 undantas 4
32916 under 916
32917 underarmen 1
32918 underbar 4
32919 underbara 2
32920 underbart 5
32921 underblåsa 1
32922 underblåser 3
32923 underbygga 1
32924 underbyggda 2
32925 undercover-verksamhet 1
32926 underfinansierade 1
32927 underformulär 1
32928 underfund 3
32929 underförstådd 1
32930 underförstås 1
32931 underförstått 1
32932 undergräva 5
32933 undergrävas 3
32934 undergräver 3
32935 undergrävs 1
32936 undergång 1
32937 undergår 1
32938 underhandsrapport 1
32939 underhus 1
32940 underhuset 4
32941 underhåll 5
32942 underhåller 1
32943 underhållet 2
32944 underhållna 1
32945 underhållningsbranschen 1
32946 underhålls 1
32947 underjordiska 4
32948 underkasta 4
32949 underkastad 1
32950 underkastas 2
32951 underkastat 1
32952 underkastelse 1
32953 underkastelsen 1
32954 underkategori 2
32955 underlag 8
32956 underlaget 1
32957 underleverantörer 4
32958 underleverantörsområdet 1
32959 underlig 1
32960 underliga 3
32961 underliggande 9
32962 underligt 2
32963 underläge 2
32964 underlägset 1
32965 underlägsna 3
32966 underläpp 1
32967 underlätta 37
32968 underlättar 10
32969 underlättats 1
32970 underlåtande 1
32971 underlåtenhet 3
32972 underlåtenheten 1
32973 underlåter 4
32974 underlåtit 2
32975 undermappar 1
32976 undermeningen 1
32977 underminera 2
32978 underminerar 1
32979 undermineras 1
32980 undermålig 1
32981 undermåliga 1
32982 undernärda 1
32983 underordnad 2
32984 underordnade 2
32985 underordnande 1
32986 underordnas 4
32987 underordnat 1
32988 underprivilegierade 1
32989 underprogram 1
32990 underpunkt 4
32991 underrapporter 2
32992 underrepresentation 3
32993 underrepresentationen 1
32994 underrepresenterade 5
32995 underrätta 1
32996 underrättas 1
32997 underrättat 1
32998 underrättelsetjänst 1
32999 underrättelsetjänsten 1
33000 underrättelsetjänster 1
33001 underrättelsetjänsternas 1
33002 underrättelseverksamheten 1
33003 underskatta 2
33004 underskattad 1
33005 underskattade 1
33006 underskattas 2
33007 underskattat 1
33008 underskott 21
33009 underskotten 6
33010 underskottet 16
33011 underskrider 1
33012 underskrift 2
33013 underskrifter 1
33014 understiger 1
33015 understruken 1
33016 understrukit 3
33017 understrukits 2
33018 understrukna 1
33019 understryka 46
33020 understrykas 5
33021 understryker 11
33022 understryks 7
33023 underströk 7
33024 underströks 1
33025 underström 1
33026 underställa 1
33027 underställas 4
33028 underställd 3
33029 underställda 2
33030 underställs 2
33031 underställt 2
33032 underställts 1
33033 understå 1
33034 understöd 1
33035 understöddes 1
33036 understöder 2
33037 understödja 3
33038 understödjande 1
33039 understödjas 3
33040 understöds 1
33041 understödspolitik 1
33042 undersysselsättningens 1
33043 undersåte 1
33044 undersöka 35
33045 undersökande 2
33046 undersökas 10
33047 undersöker 4
33048 undersökning 22
33049 undersökningar 20
33050 undersökningarna 3
33051 undersökningarnas 1
33052 undersökningen 7
33053 undersökningsgrupp 1
33054 undersökningskommission 1
33055 undersökningskommitté 1
33056 undersökningskommittén 1
33057 undersökningsmakt 1
33058 undersökningsmekanismer 1
33059 undersökningsprocess 2
33060 undersökningssystem 1
33061 undersökt 6
33062 undersökta 2
33063 undersökte 1
33064 underteckna 6
33065 undertecknad 1
33066 undertecknade 2
33067 undertecknades 9
33068 undertecknande 1
33069 undertecknandet 1
33070 undertecknar 5
33071 undertecknarna 1
33072 undertecknas 3
33073 undertecknat 17
33074 undertecknats 4
33075 undertrycka 4
33076 undertrycker 2
33077 undertryckta 1
33078 underutnyttjande 1
33079 underutvecklad 3
33080 underutvecklade 3
33081 underutvecklat 1
33082 underutveckling 2
33083 underutvecklingen 2
33084 undervattensfloder 1
33085 undervattenssamling 1
33086 undervegetationen 1
33087 underverk 1
33088 undervisa 1
33089 undervisade 1
33090 undervisat 1
33091 undervisning 3
33092 undervisningen 2
33093 undervärdera 1
33094 undfallande 1
33095 undgick 1
33096 undgå 3
33097 undgår 3
33098 undgått 3
33099 undkomma 2
33100 undkommer 2
33101 undkommit 2
33102 undlåtit 1
33103 undra 5
33104 undrade 11
33105 undran 4
33106 undrande 2
33107 undrar 41
33108 undsluppit 1
33109 undsätta 1
33110 undvik 1
33111 undvika 90
33112 undvikas 8
33113 undviker 8
33114 undvikit 4
33115 undvikits 1
33116 undviks 2
33117 ung 23
33118 ung. 1
33119 unga 40
33120 ungdom 3
33121 ungdomar 23
33122 ungdomarna 3
33123 ungdomarnas 1
33124 ungdomen 2
33125 ungdomlig 1
33126 ungdoms- 3
33127 ungdomsarbetslöshet 2
33128 ungdomsarbetslösheten 1
33129 ungdomsbrottslighet 3
33130 ungdomsfrågor 3
33131 unge 13
33132 ungefär 21
33133 ungefärliga 1
33134 ungerska 1
33135 ungfisken 1
33136 ungkarl 1
33137 ungkarlarna 1
33138 ungrare 1
33139 ungt 1
33140 uniform 2
33141 uniformer 1
33142 uniformerade 1
33143 unik 4
33144 unika 12
33145 unikt 6
33146 unilaterala 2
33147 unilateralt 3
33148 union 60
33149 unionen 854
33150 unionen-Afrika 2
33151 unionen-Kina 1
33152 unionens 406
33153 unions 1
33154 unions- 1
33155 unionsfördrag 1
33156 unionsfördraget 1
33157 unionsmedborgare 2
33158 unionsmedborgarna 1
33159 unionsmedborgarnas 2
33160 unionsmedlemmar 1
33161 unionsnivå 6
33162 unionssammanhang 1
33163 universalitet 1
33164 universaliteten 1
33165 universalmedel 1
33166 universell 3
33167 universella 10
33168 universitet 2
33169 universiteten 1
33170 universitetet 4
33171 universitetsmiljöerna 1
33172 universum 1
33173 universums 2
33174 unna 1
33175 uns 1
33176 unset 1
33177 upp 837
33178 upp-land 1
33179 uppassade 1
33180 uppassare 1
33181 uppbackning 1
33182 uppbjuda 1
33183 uppblandad 1
33184 uppblandning 1
33185 uppblötta 1
33186 uppborstat 1
33187 uppbringa 1
33188 uppbringar 2
33189 uppbringas 2
33190 uppbromsningen 1
33191 uppbrottsstämning 1
33192 uppburits 1
33193 uppbyggande 1
33194 uppbyggandet 1
33195 uppbyggd 1
33196 uppbyggnad 5
33197 uppbyggnaden 16
33198 uppbyggnadsplatserna 1
33199 uppbyggt 4
33200 uppbär 1
33201 uppbära 2
33202 uppbåda 2
33203 uppdatera 6
33204 uppdaterad 1
33205 uppdateras 1
33206 uppdatering 1
33207 uppdelad 1
33208 uppdelade 1
33209 uppdelat 4
33210 uppdelning 4
33211 uppdelningen 4
33212 uppdrag 41
33213 uppdragen 1
33214 uppdraget 5
33215 uppdragna 1
33216 uppdrog 1
33217 uppdykandet 1
33218 uppe 16
33219 uppehälle 2
33220 uppehåll 2
33221 uppehålla 12
33222 uppehåller 4
33223 uppehållet 1
33224 uppehållit 1
33225 uppehållstillstånd 5
33226 uppehållstillståndet 2
33227 uppehållstillståndets 1
33228 uppehållsvillkor 1
33229 uppenbar 6
33230 uppenbara 6
33231 uppenbarar 1
33232 uppenbarelse 2
33233 uppenbarelse-kvalitet 1
33234 uppenbarligen 31
33235 uppenbart 69
33236 uppfanns 1
33237 uppfatta 2
33238 uppfattade 4
33239 uppfattar 20
33240 uppfattas 6
33241 uppfattat 3
33242 uppfattbart 1
33243 uppfattning 71
33244 uppfattningar 10
33245 uppfattningen 13
33246 uppfinna 3
33247 uppfinning 2
33248 uppfinningarnas 1
33249 uppfostrades 1
33250 uppfostran 2
33251 uppfostrat 1
33252 uppfriskande 1
33253 uppfylla 60
33254 uppfyllandet 6
33255 uppfyllas 11
33256 uppfylld 2
33257 uppfyllda 4
33258 uppfyllde 3
33259 uppfylldes 2
33260 uppfyller 37
33261 uppfylls 8
33262 uppfyllt 1
33263 uppfyllts 5
33264 uppfångade 1
33265 uppfödning 1
33266 uppföljas 1
33267 uppföljning 15
33268 uppföljningen 6
33269 uppföljningsfråga 1
33270 uppföljningskommittén 2
33271 uppföljningsrapporten 1
33272 uppföljningsregler 1
33273 uppför 13
33274 uppföra 4
33275 uppförande 5
33276 uppförandekod 6
33277 uppförandekoden 3
33278 uppförandekoder 2
33279 uppförandekoderna 1
33280 uppföranderegler 2
33281 uppförandereglerna 1
33282 uppförandet 3
33283 uppförde 2
33284 uppförs 1
33285 uppförstorad 1
33286 uppfört 1
33287 uppgavs 1
33288 uppger 1
33289 uppges 1
33290 uppgick 5
33291 uppgift 98
33292 uppgiften 9
33293 uppgifter 130
33294 uppgifterna 27
33295 uppgifternas 1
33296 uppgiftsfördelning 1
33297 uppgiftslämnare 1
33298 uppgiftsmängd 1
33299 uppgivande 1
33300 uppgradera 1
33301 uppgå 3
33302 uppgående 1
33303 uppgång 3
33304 uppgången 1
33305 uppgår 14
33306 uppgörelse 3
33307 uppgörelsen 2
33308 uppgörelser 2
33309 uppgörelserna 2
33310 upphandling 2
33311 upphetsad 1
33312 upphetsade 1
33313 upphetsande 1
33314 upphetsat 1
33315 upphetsning 1
33316 upphettat 1
33317 upphov 33
33318 upphovet 1
33319 upphovskällan 1
33320 upphovsman 4
33321 upphovsmannen 2
33322 upphovsmän 2
33323 upphovsmännen 4
33324 upphovsmännens 1
33325 upphovsrätt 11
33326 upphovsrätten 4
33327 upphovsrättsavgift 1
33328 upphovsrättsliga 1
33329 upphovsrättsligt 1
33330 upphovsrättsreglering 1
33331 upphängd 1
33332 upphängda 1
33333 upphäva 8
33334 upphävande 2
33335 upphävandet 3
33336 upphävas 5
33337 upphävdes 1
33338 upphävs 2
33339 upphöja 1
33340 upphöjd 1
33341 upphöjda 2
33342 upphöjs 1
33343 upphör 7
33344 upphöra 14
33345 upphörandet 1
33346 upphörde 5
33347 upphört 7
33348 uppifrån 2
33349 uppkallad 1
33350 uppklädd 1
33351 uppkomma 2
33352 uppkommer 8
33353 uppkommit 5
33354 uppkomsten 1
33355 upplagan 1
33356 uppleva 15
33357 upplevde 5
33358 upplevelse 4
33359 upplevelser 1
33360 upplevelses 1
33361 upplever 14
33362 upplevs 2
33363 upplevt 6
33364 upplyftande 1
33365 upplysa 7
33366 upplyses 1
33367 upplysning 6
33368 upplysningar 5
33369 upplyst 7
33370 upplysta 4
33371 upplyste 2
33372 upplysts 1
33373 upplåsta 1
33374 upplösa 1
33375 upplöses 1
33376 upplösning 7
33377 upplösta 1
33378 upplöstes 2
33379 uppmana 28
33380 uppmanade 5
33381 uppmanades 1
33382 uppmanar 69
33383 uppmanas 12
33384 uppmanat 3
33385 uppmaning 12
33386 uppmaningar 3
33387 uppmaningen 2
33388 uppmaningsskrivelse 1
33389 uppmjukning 3
33390 uppmjukningen 2
33391 uppmuntra 37
33392 uppmuntrad 1
33393 uppmuntran 5
33394 uppmuntrande 9
33395 uppmuntrar 18
33396 uppmuntras 13
33397 uppmuntrat 2
33398 uppmuntrats 1
33399 uppmärksam 5
33400 uppmärksamhet 80
33401 uppmärksamheten 17
33402 uppmärksamma 23
33403 uppmärksammade 2
33404 uppmärksammar 4
33405 uppmärksammare 1
33406 uppmärksammas 7
33407 uppmärksammat 2
33408 uppmärksammats 1
33409 uppmärksamt 12
33410 uppmätta 1
33411 uppmättes 1
33412 uppnå 139
33413 uppnåbara 1
33414 uppnådda 6
33415 uppnådde 3
33416 uppnåddes 2
33417 uppnåeligt 1
33418 uppnår 21
33419 uppnås 36
33420 uppnått 20
33421 uppnåtts 17
33422 uppochner 1
33423 uppochnervända 1
33424 uppoffrande 1
33425 uppoffrat 1
33426 uppoffring 1
33427 uppoffringar 2
33428 upprensningar 1
33429 upprensningen 1
33430 upprepa 38
33431 upprepade 29
33432 upprepades 1
33433 upprepandets 1
33434 upprepar 41
33435 upprepas 15
33436 upprepat 4
33437 upprepats 3
33438 upprepning 2
33439 uppriktig 1
33440 uppriktiga 2
33441 uppriktighet 1
33442 uppriktigt 15
33443 uppritade 1
33444 upprivande 1
33445 upprop 2
33446 uppror 1
33447 upproriska 1
33448 upprusta 1
33449 uppryckning 1
33450 uppräknade 1
33451 uppräkning 2
33452 upprätta 29
33453 upprättade 2
33454 upprättades 1
33455 upprättande 4
33456 upprättandet 10
33457 upprättar 14
33458 upprättas 6
33459 upprättat 9
33460 upprättats 3
33461 upprättelse 1
33462 upprätthålla 20
33463 upprätthållande 1
33464 upprätthållandet 4
33465 upprätthållas 2
33466 upprätthåller 3
33467 upprätthållit 1
33468 upprätthålls 3
33469 uppröjningsarbetet 1
33470 uppröra 1
33471 upprörande 5
33472 uppröras 1
33473 upprörd 2
33474 upprörda 2
33475 upprördhet 1
33476 uppsamling 3
33477 uppsamlingen 1
33478 uppsamlingscentrum 1
33479 uppsamlingsplatser 2
33480 uppsamlingsplatserna 1
33481 uppsatt 4
33482 uppsatta 4
33483 uppseendeväckande 3
33484 uppsjö 1
33485 uppskakade 1
33486 uppskatta 9
33487 uppskattad 1
33488 uppskattade 4
33489 uppskattande 2
33490 uppskattar 22
33491 uppskattas 3
33492 uppskattat 1
33493 uppskattning 16
33494 uppskattningar 2
33495 uppskattningsvis 1
33496 uppskjuta 2
33497 uppskjutande 3
33498 uppskjutas 2
33499 uppskjuten 1
33500 uppskjuter 1
33501 uppskov 1
33502 uppskovet 1
33503 uppskruvade 3
33504 uppslagen 1
33505 uppslitsade 1
33506 uppsluppna 1
33507 uppsluppnaste 1
33508 uppslutning 1
33509 uppspaltning 1
33510 uppspelt 1
33511 uppsplittring 1
33512 uppspärrade 1
33513 uppspårandet 1
33514 uppspårningsfasen 1
33515 uppstaplade 1
33516 uppstod 8
33517 uppstoppade 1
33518 uppsträckta 1
33519 uppströms 5
33520 uppställa 2
33521 uppställandet 1
33522 uppställas 1
33523 uppställda 5
33524 uppställer 1
33525 uppställning 1
33526 uppställningsspår 1
33527 uppstå 17
33528 uppståndelse 1
33529 uppståndelsen 1
33530 uppstår 47
33531 uppstått 19
33532 uppsving 5
33533 uppsyn 1
33534 uppsägning 1
33535 uppsägningar 11
33536 uppsägningsbesked 1
33537 uppsägningsbeskedet 1
33538 uppsättning 5
33539 upptagen 5
33540 upptaget 4
33541 upptagetton 1
33542 upptagit 1
33543 upptagits 1
33544 upptagna 2
33545 upptagningsområde 1
33546 upptar 3
33547 upptas 3
33548 upptrappningen 1
33549 uppträda 2
33550 uppträdande 9
33551 uppträdde 1
33552 uppträder 8
33553 uppträtt 1
33554 upptäcka 7
33555 upptäckas 1
33556 upptäcker 6
33557 upptäcks 3
33558 upptäckt 7
33559 upptäckte 17
33560 upptäckten 3
33561 upptäcktes 3
33562 upptäckts 5
33563 upptäcktsfärdernas 1
33564 uppvaknad 1
33565 uppviglande 1
33566 uppvisa 5
33567 uppvisade 1
33568 uppvisar 11
33569 uppvisas 1
33570 uppvisat 4
33571 uppvisning 1
33572 uppväga 3
33573 uppväger 1
33574 uppvända 1
33575 uppvärdera 1
33576 uppvärderar 2
33577 uppvärdering 2
33578 uppäten 1
33579 uppåt 8
33580 uppåtseende 1
33581 ur 157
33582 uran 8
33583 uranium 2
33584 uranvapen 4
33585 urartad 1
33586 urartade 1
33587 urartande 1
33588 urartar 1
33589 urban 3
33590 urbana 4
33591 urbanisering 1
33592 urbaniseringen 2
33593 urgamla 1
33594 urgammal 1
33595 urholka 3
33596 urholkar 1
33597 urholkas 4
33598 urholkat 1
33599 urholkningen 1
33600 urminnes 1
33601 urringning 1
33602 ursinnig 1
33603 urskilja 6
33604 urskiljas 1
33605 urskiljer 3
33606 urskillningslöst 1
33607 urskogar 1
33608 urskuldande 1
33609 ursprung 25
33610 ursprunget 6
33611 ursprungliga 51
33612 ursprungligen 9
33613 ursprungsbefolkning 1
33614 ursprungsbefolkningar 4
33615 ursprungsbestämmelser 1
33616 ursprungsfrågor 1
33617 ursprungsintyg 1
33618 ursprungskick 1
33619 ursprungsland 2
33620 ursprungslandet 1
33621 ursprungsländer 1
33622 ursprungsländerna 3
33623 ursprungsmärkning 1
33624 ursprungsregionerna 1
33625 ursprungsregler 2
33626 ursprungsreglerna 1
33627 ursprungsversionen 1
33628 urspårning 1
33629 ursäkt 21
33630 ursäkta 9
33631 ursäktade 1
33632 ursäktande 2
33633 ursäktar 1
33634 ursäkten 2
33635 ursäkter 4
33636 urtider 1
33637 urval 5
33638 urvalet 5
33639 urvalsfråga 2
33640 urvalsfrågan 1
33641 urvalskommittéerna 1
33642 urvalskriterier 2
33643 urvalskriterierna 2
33644 urvattna 2
33645 urvattnade 1
33646 urvattnar 2
33647 urvattnas 3
33648 urvattnat 1
33649 urvattning 3
33650 uråldriga 1
33651 uråldrigare 1
33652 ut 536
33653 ut-och-invändningsteknik 1
33654 utan 953
33655 utanför 107
33656 utanförskap 3
33657 utanpå 1
33658 utantill 1
33659 utarbeta 43
33660 utarbetade 6
33661 utarbetades 3
33662 utarbetande 1
33663 utarbetandet 19
33664 utarbetar 9
33665 utarbetas 9
33666 utarbetat 9
33667 utarbetats 6
33668 utarmade 5
33669 utarmar 1
33670 utarmas 1
33671 utarmat 6
33672 utarmningen 1
33673 utbasunerade 1
33674 utbetalade 3
33675 utbetalades 1
33676 utbetalas 1
33677 utbetalning 3
33678 utbetalningar 1
33679 utbetalningarna 1
33680 utbetalningen 3
33681 utbilda 4
33682 utbildade 4
33683 utbildar 2
33684 utbildas 4
33685 utbildats 1
33686 utbildning 65
33687 utbildningar 2
33688 utbildningen 9
33689 utbildningens 1
33690 utbildnings- 5
33691 utbildningscentra 1
33692 utbildningscentren 1
33693 utbildningsinsatser 1
33694 utbildningsinstitutioner 2
33695 utbildningskostnader 2
33696 utbildningsministern 1
33697 utbildningsmoment 1
33698 utbildningsmöjligheter 1
33699 utbildningsnivå 3
33700 utbildningsnivån 1
33701 utbildningsoffensiv 1
33702 utbildningsområdet 1
33703 utbildningspolitiken 2
33704 utbildningspolitisk 2
33705 utbildningspraktik 1
33706 utbildningsprogram 2
33707 utbildningsprojekt 1
33708 utbildningssamhälle 1
33709 utbildningsstrukturer 1
33710 utbildningssystem 1
33711 utbildningssystemens 1
33712 utbildningssystemet 1
33713 utbildningsåtgärder 1
33714 utblottade 1
33715 utbrast 1
33716 utbredd 3
33717 utbredda 1
33718 utbredning 6
33719 utbredningen 1
33720 utbrister 1
33721 utbrott 3
33722 utbrottet 1
33723 utbrutit 1
33724 utbrytarstyrkor 1
33725 utbud 6
33726 utbudet 2
33727 utbudsinriktad 1
33728 utbyggd 1
33729 utbyggnad 4
33730 utbyggnaden 2
33731 utbyggt 1
33732 utbyta 5
33733 utbyte 30
33734 utbyten 1
33735 utbyter 2
33736 utbytesprincipen 1
33737 utbytesprojekt 2
33738 utbytet 7
33739 utbytte 2
33740 utbärningar 1
33741 utdata 1
33742 utdela 1
33743 utdelad 1
33744 utdelar 1
33745 utdelas 2
33746 utdelning 3
33747 utdelningen 2
33748 utdrag 1
33749 utdragen 2
33750 utdragna 2
33751 utdömda 1
33752 utdömer 2
33753 ute 37
33754 uteblivit 1
33755 utedasset 1
33756 utefter 1
33757 utelämna 1
33758 utelämnade 1
33759 utelämnas 4
33760 utesluta 6
33761 uteslutande 15
33762 uteslutas 2
33763 utesluten 1
33764 utesluter 7
33765 uteslutet 2
33766 uteslutits 1
33767 uteslutna 1
33768 uteslutning 6
33769 utesluts 1
33770 uteslöt 2
33771 utestänga 1
33772 utestängas 4
33773 utestängda 1
33774 utestängning 2
33775 utestängs 1
33776 utestängt 1
33777 utestängts 1
33778 utfall 1
33779 utfallet 1
33780 utfarten 1
33781 utfasning 3
33782 utfasningen 4
33783 utfiskning 1
33784 utflaggningsländer 1
33785 utflykter 2
33786 utflyttade 1
33787 utflyttningen 1
33788 utflyttningsbidrag 1
33789 utfodrat 1
33790 utforma 25
33791 utformad 3
33792 utformade 9
33793 utformades 1
33794 utformandet 3
33795 utformar 6
33796 utformas 13
33797 utformat 4
33798 utformats 1
33799 utformning 21
33800 utformningar 1
33801 utformningen 21
33802 utformningsmässiga 1
33803 utforska 2
33804 utforskas 1
33805 utfrågning 9
33806 utfrågningar 1
33807 utfrågningarna 1
33808 utfrågningen 4
33809 utfärda 8
33810 utfärdades 1
33811 utfärdande 4
33812 utfärdandet 2
33813 utfärdar 1
33814 utfärdas 1
33815 utfärdat 3
33816 utfärdats 1
33817 utfästelser 2
33818 utför 13
33819 utföra 29
33820 utförande 2
33821 utföras 2
33822 utförd 1
33823 utförda 2
33824 utförde 2
33825 utfördes 2
33826 utförlig 2
33827 utförliga 2
33828 utförligare 1
33829 utförligen 1
33830 utförligt 2
33831 utförs 8
33832 utfört 13
33833 utförts 6
33834 utgallring 4
33835 utgallringen 1
33836 utgavs 1
33837 utgick 3
33838 utgifter 27
33839 utgifterna 11
33840 utgifts 1
33841 utgiftsmål 1
33842 utgiftsområde 11
33843 utgiftsområden 1
33844 utgiftsområdet 1
33845 utgiftspolitik 1
33846 utgiftsprioriteringar 1
33847 utgiftsprogram 1
33848 utgiftssektorer 1
33849 utgiftstak 1
33850 utgivare 1
33851 utgivit 1
33852 utgivna 2
33853 utgjorde 10
33854 utgjordes 1
33855 utgjort 3
33856 utgrävningen 1
33857 utgå 11
33858 utgång 4
33859 utgången 9
33860 utgångsförslag 1
33861 utgångsläge 1
33862 utgångspunkt 22
33863 utgångspunkten 5
33864 utgångspunkter 4
33865 utgår 25
33866 utgått 4
33867 utgåva 1
33868 utgåvor 1
33869 utgör 135
33870 utgöra 34
33871 utgörs 8
33872 utgör­ 1
33873 uthuset 1
33874 uthyrning 5
33875 uthärda 1
33876 uthärdliga 1
33877 uthållighet 2
33878 utifrån 48
33879 utjämna 4
33880 utjämningen 1
33881 utjämningsfond 1
33882 utkanten 5
33883 utkast 13
33884 utkasten 1
33885 utkastet 10
33886 utkik 1
33887 utkom 1
33888 utkomst 3
33889 utkonkurrerade 1
33890 utkräva 1
33891 utkrävandet 1
33892 utkräver 2
33893 utkämpa 2
33894 utkämpar 1
33895 utlandet 4
33896 utlandsplacerade 2
33897 utlandsplacering 1
33898 utloppet 1
33899 utlovade 7
33900 utlovar 1
33901 utlovat 3
33902 utlovats 1
33903 utlyst 2
33904 utlägg 1
33905 utläggningar 1
33906 utlämna 1
33907 utlämnad 1
33908 utlämnats 1
33909 utlämning 1
33910 utländsk 2
33911 utländska 12
33912 utlänningslagarna 1
33913 utlänningslagen 2
33914 utläsa 1
33915 utlåning 2
33916 utlåtande 1
33917 utlåtanden 1
33918 utlåtandet 1
33919 utlösa 1
33920 utlösande 1
33921 utlöst 1
33922 utlöste 1
33923 utlöstes 1
33924 utmana 3
33925 utmanande 3
33926 utmanas 1
33927 utmaning 31
33928 utmaningar 37
33929 utmaningarna 7
33930 utmaningen 15
33931 utmattad 1
33932 utmattning 1
33933 utmed 4
33934 utmynnar 1
33935 utmynnat 1
33936 utmärkande 1
33937 utmärker 3
33938 utmärks 2
33939 utmärkt 48
33940 utmärkta 40
33941 utnyttja 56
33942 utnyttjade 2
33943 utnyttjades 3
33944 utnyttjande 14
33945 utnyttjandet 7
33946 utnyttjar 11
33947 utnyttjas 19
33948 utnyttjat 5
33949 utnyttjats 1
33950 utnämna 3
33951 utnämnandet 1
33952 utnämndes 1
33953 utnämner 1
33954 utnämning 1
33955 utnämningen 1
33956 utnämnt 1
33957 utnämnts 2
33958 utom 17
33959 utomeuropeiska 6
33960 utomeuropeiskt 1
33961 utomhus 1
33962 utomlands 2
33963 utomordentlig 1
33964 utomordentliga 3
33965 utomordentligt 16
33966 utomstående 6
33967 utopier 1
33968 utopiskt 1
33969 utpeka 1
33970 utpekar 1
33971 utpekas 1
33972 utplacerad 1
33973 utplacerade 2
33974 utplacerades 1
33975 utplacering 2
33976 utplåna 4
33977 utplånade 1
33978 utplånande 1
33979 utplånar 1
33980 utplånat 1
33981 utplåning 3
33982 utpressning 3
33983 utpräglad 1
33984 utpräglade 1
33985 utrangeras 1
33986 utreda 3
33987 utredande 2
33988 utredd 1
33989 utredning 4
33990 utredningar 5
33991 utredningarna 1
33992 utredningsarbetet 1
33993 utredningsbyråer 1
33994 utredningshäktning 1
33995 utredningstekniska 1
33996 utredningsverksamhet 1
33997 utreds 1
33998 utrikes 3
33999 utrikes- 21
34000 utrikesdepartementet 3
34001 utrikesenhet 1
34002 utrikesfrågor 13
34003 utrikesförbindelser 2
34004 utrikeshandel 5
34005 utrikeshandelspolitikerna 1
34006 utrikeskorrespondenter 1
34007 utrikesminister 4
34008 utrikesministeriernas 1
34009 utrikesministern 7
34010 utrikesministrarna 2
34011 utrikesnivå 1
34012 utrikespolitik 12
34013 utrikespolitiken 15
34014 utrikespolitisk 1
34015 utrikespolitiska 4
34016 utropa 1
34017 utropar 1
34018 utropas 2
34019 utrota 16
34020 utrotad 1
34021 utrotas 2
34022 utrotning 2
34023 utrotningar 1
34024 utrotningen 2
34025 utrotningshotade 1
34026 utrotningsstrategier 1
34027 utrotningsåtgärder 1
34028 utrullad 1
34029 utrustad 1
34030 utrustade 1
34031 utrustar 2
34032 utrustas 2
34033 utrustning 8
34034 utrustningar 1
34035 utrustningen 2
34036 utrymme 24
34037 utrymmet 2
34038 uträtta 6
34039 uträttar 1
34040 uträttat 2
34041 utröna 3
34042 utsatt 5
34043 utsatta 10
34044 utsattes 1
34045 utsatthet 1
34046 utsatts 3
34047 utse 4
34048 utsedd 1
34049 utsedda 2
34050 utseende 13
34051 utseendet 1
34052 utser 2
34053 utses 3
34054 utsett 2
34055 utsetts 1
34056 utsikt 6
34057 utsikten 3
34058 utsikter 4
34059 utsikterna 5
34060 utsirade 1
34061 utskott 60
34062 utskotten 7
34063 utskottet 293
34064 utskottets 16
34065 utskotts 3
34066 utskottsbehandlingen 5
34067 utskottsdebatten 1
34068 utskottsförhandlingen 1
34069 utskottsrummen 1
34070 utskottssammanträdet 1
34071 utskottssekretariatet 1
34072 utslag 3
34073 utslagen 1
34074 utslagna 4
34075 utslagning 20
34076 utslagningen 6
34077 utslagningens 1
34078 utslagningsmekanismer 1
34079 utslagningspolitik 1
34080 utslungade 1
34081 utsläpp 15
34082 utsläppen 11
34083 utsläppet 5
34084 utsläppsnivåer 1
34085 utsläppsrätter 1
34086 utslätning 1
34087 utspelad 1
34088 utspelade 2
34089 utspridd 1
34090 utspridda 3
34091 utspridning 1
34092 utspärrade 1
34093 utstationera 1
34094 utstationerad 1
34095 utstationerade 1
34096 utstationering 7
34097 utstationeringssituationen 1
34098 utsträcka 1
34099 utsträckas 2
34100 utsträckning 69
34101 utsträckningen 1
34102 utsträcks 1
34103 utsträckt 1
34104 utsträckta 1
34105 utstrålade 1
34106 utstrålar 1
34107 utströdda 1
34108 utstuderad 2
34109 utställandet 1
34110 utställda 1
34111 utställningar 4
34112 utställningsföremål 1
34113 utställt 1
34114 utstå 5
34115 utstående 2
34116 utstår 1
34117 utstått 2
34118 utstötta 3
34119 utsugare 2
34120 utsugning 1
34121 utsvulten 1
34122 utsäde 4
34123 utsända 1
34124 utsätta 6
34125 utsättas 5
34126 utsätter 1
34127 utsättningsdirektivet 1
34128 utsätts 11
34129 utsågs 3
34130 utsålda 1
34131 utsökta 1
34132 utsöndrade 1
34133 uttag 1
34134 uttagningsprov 1
34135 uttala 39
34136 uttalad 3
34137 uttalade 17
34138 uttalades 3
34139 uttalande 89
34140 uttalanden 47
34141 uttalandena 4
34142 uttalandet 10
34143 uttalar 17
34144 uttalas 4
34145 uttalat 17
34146 uttaxeraren 1
34147 uttjänta 25
34148 uttolkare 1
34149 uttolkarna 1
34150 uttorkning 2
34151 uttrar 1
34152 uttryck 67
34153 uttrycka 48
34154 uttryckas 2
34155 uttrycker 13
34156 uttrycket 9
34157 uttrycklig 2
34158 uttryckliga 3
34159 uttryckligen 20
34160 uttryckligt 1
34161 uttrycks 13
34162 uttrycksfull 1
34163 uttryckslös 1
34164 uttryckt 16
34165 uttryckta 2
34166 uttryckte 21
34167 uttrycktes 3
34168 uttryckts 4
34169 utträda 1
34170 utträde 1
34171 uttänkt 1
34172 uttänkta 1
34173 uttömd 1
34174 uttömda 1
34175 uttömmande 6
34176 uttömt 1
34177 utvald 1
34178 utvalda 2
34179 utvandring 2
34180 utveckla 77
34181 utvecklad 4
34182 utvecklade 33
34183 utvecklades 2
34184 utvecklande 2
34185 utvecklandet 3
34186 utvecklar 8
34187 utvecklare 3
34188 utvecklaren 4
34189 utvecklas 59
34190 utvecklat 9
34191 utvecklats 13
34192 utveckling 285
34193 utvecklingar 1
34194 utvecklingen 169
34195 utvecklingens 2
34196 utvecklings- 9
34197 utvecklingsaktörer 1
34198 utvecklingsarbete 1
34199 utvecklingsaspekterna 1
34200 utvecklingsbistånd 7
34201 utvecklingsbiståndet 1
34202 utvecklingsbiståndsprogram 1
34203 utvecklingsbudget 1
34204 utvecklingscentrum 1
34205 utvecklingscentrumet 1
34206 utvecklingsfas 2
34207 utvecklingsfond 1
34208 utvecklingsfonden 15
34209 utvecklingsfondens 1
34210 utvecklingsfonder 1
34211 utvecklingsfrämjande 1
34212 utvecklingsfråga 2
34213 utvecklingsfrågan 1
34214 utvecklingsfrågor 3
34215 utvecklingsfunktioner 1
34216 utvecklingsfunktionerna 1
34217 utvecklingsförmåga 1
34218 utvecklingshjälp 1
34219 utvecklingshjälpen 1
34220 utvecklingsinitiativ 1
34221 utvecklingsinsatser 1
34222 utvecklingsinstrument 1
34223 utvecklingskonferens 1
34224 utvecklingsland 1
34225 utvecklingsländer 15
34226 utvecklingsländerna 42
34227 utvecklingsländernas 7
34228 utvecklingsmetod 1
34229 utvecklingsminister 1
34230 utvecklingsmodell 2
34231 utvecklingsmässigt 1
34232 utvecklingsmål 1
34233 utvecklingsmålen 3
34234 utvecklingsmöjligheter 1
34235 utvecklingsmöjligheterna 1
34236 utvecklingsmönster 1
34237 utvecklingsnationerna 2
34238 utvecklingsnivå 1
34239 utvecklingsnivåer 2
34240 utvecklingsområde 1
34241 utvecklingsområden 1
34242 utvecklingsområdet 3
34243 utvecklingspartner 2
34244 utvecklingspartnerskap 4
34245 utvecklingspartnerskapen 1
34246 utvecklingspartnerskapens 1
34247 utvecklingsperspektivet 1
34248 utvecklingsplan 1
34249 utvecklingsplanerna 1
34250 utvecklingspolicy 1
34251 utvecklingspolitik 14
34252 utvecklingspolitiken 36
34253 utvecklingspotential 1
34254 utvecklingsprioriteringar 1
34255 utvecklingsprioriteringarna 1
34256 utvecklingsprocess 2
34257 utvecklingsprocessen 1
34258 utvecklingsprogram 4
34259 utvecklingsprogrammen 6
34260 utvecklingsprojekt 2
34261 utvecklingsprojekten 1
34262 utvecklingsprojekts 1
34263 utvecklingsredskapet 1
34264 utvecklingssamarbete 9
34265 utvecklingssamarbetesaspekten 1
34266 utvecklingssamarbetet 5
34267 utvecklingssamhället 1
34268 utvecklingsstadiet 2
34269 utvecklingssteg 1
34270 utvecklingsstrategi 1
34271 utvecklingsstrategier 3
34272 utvecklingsstrategierna 1
34273 utvecklingsstöd 6
34274 utvecklingsstödet 1
34275 utvecklingstakten 1
34276 utvecklingstjänstemän 1
34277 utvecklingstjänsterna 1
34278 utvecklingsväg 1
34279 utvecklingsändamål 1
34280 utverka 5
34281 utvidga 28
34282 utvidgad 5
34283 utvidgade 3
34284 utvidgades 1
34285 utvidgande 1
34286 utvidgar 8
34287 utvidgas 18
34288 utvidgat 3
34289 utvidgning 49
34290 utvidgningar 2
34291 utvidgningarna 1
34292 utvidgningen 99
34293 utvidgningens 4
34294 utvidgningsfrågan 1
34295 utvidgningsplanerna 1
34296 utvidgningsprocess 1
34297 utvidgningsprocessen 6
34298 utvidgningsprojektet 2
34299 utvidgningsrunda 1
34300 utvidgningsärendet 1
34301 utvinningsnivåer 1
34302 utvinns 1
34303 utvisa 3
34304 utvisade 1
34305 utvisar 1
34306 utvisning 4
34307 utväg 5
34308 utvärdera 12
34309 utvärderar 2
34310 utvärderas 6
34311 utvärderat 1
34312 utvärdering 30
34313 utvärderingar 6
34314 utvärderingarna 1
34315 utvärderingen 15
34316 utvärderingskommittéerna 1
34317 utvärderingspanelerna 1
34318 utväxlade 2
34319 utväxlandet 1
34320 utväxlat 1
34321 utväxling 2
34322 utåt 5
34323 utöka 13
34324 utökad 2
34325 utökade 1
34326 utökades 2
34327 utökande 1
34328 utökar 2
34329 utökas 4
34330 utökat 3
34331 utökning 2
34332 utöva 18
34333 utövade 1
34334 utövades 1
34335 utövande 9
34336 utövandet 2
34337 utövar 9
34338 utövas 9
34339 utövat 1
34340 utöver 24
34341 v 1
34342 va 4
34343 vaccin 10
34344 vaccination 2
34345 vaccinationsprogram 1
34346 vacciner 1
34347 vaccinera 1
34348 vaccinering 5
34349 vaccinet 1
34350 vacker 10
34351 vackert 3
34352 vackla 1
34353 vacklade 1
34354 vackra 23
34355 vackraste 2
34356 vad 771
34357 vag 2
34358 vaga 11
34359 vagabond 1
34360 vaggan 1
34361 vagnar 1
34362 vagnen 3
34363 vagt 4
34364 vajande 1
34365 vaka 2
34366 vakande 1
34367 vakanta 1
34368 vakar 2
34369 vaken 2
34370 vaket 1
34371 vakna 3
34372 vaknade 7
34373 vaknar 2
34374 vaksam 6
34375 vaksamhet 4
34376 vaksamma 10
34377 vaksammare 1
34378 vaksamt 2
34379 vakt 4
34380 vaktade 1
34381 vakter 1
34382 vaktmästarna 1
34383 vakuum 3
34384 vakuumtankar 1
34385 val 51
34386 valar 1
34387 valbarhet 1
34388 valbart 1
34389 vald 10
34390 valda 20
34391 valdagen 1
34392 valde 7
34393 valdeltagandet 7
34394 valdes 4
34395 valdistrikt 2
34396 valen 10
34397 valet 17
34398 valfläsk 1
34399 valframgång 1
34400 valframgångar 2
34401 valfrihet 1
34402 valfriheten 2
34403 valfråga 1
34404 valfusket 1
34405 valförfaranden 1
34406 validerades 1
34407 valkampanj 3
34408 valkampanjen 2
34409 valkampanjerna 1
34410 valkrets 6
34411 valkretsar 1
34412 valkretsen 1
34413 vallfärd 1
34414 vallfärdsstav 1
34415 vallistorna 2
34416 vallokalerna 1
34417 valman 1
34418 valmässiga 1
34419 valmöjligheter 2
34420 valnötsträden 1
34421 valobservation 1
34422 valobservatörer 1
34423 valområden 1
34424 valperioden 1
34425 valresultaten 1
34426 valresultatet 2
34427 valrörelse 1
34428 valrörelsen 1
34429 valsedlar 1
34430 valseger 1
34431 valt 21
34432 valtaktiska 1
34433 valtider 2
34434 valts 9
34435 valuation 1
34436 valuta 18
34437 valutafonden 4
34438 valutafondens 1
34439 valutafrågor 27
34440 valutaförfalskare 1
34441 valutaförfalskning 3
34442 valutaförfalskningar 1
34443 valutaförfalskningen 1
34444 valutaförfalskningsbrott 1
34445 valutan 21
34446 valutans 4
34447 valutapolitikens 1
34448 valutarisker 1
34449 valutaspekulationen 2
34450 valutaunionen 3
34451 valutaunionens 1
34452 valutor 5
34453 valutorna 3
34454 valv 2
34455 valven 1
34456 valörer 1
34457 valövervakningen 1
34458 vampyr 1
34459 van 38
34460 vana 4
34461 vandra 6
34462 vandrade 7
34463 vandrande 1
34464 vandrare 1
34465 vandringar 2
34466 vanhedra 1
34467 vanhedrande 2
34468 vanlig 11
34469 vanliga 23
34470 vanligare 5
34471 vanligaste 3
34472 vanligen 2
34473 vanligt 15
34474 vanligtvis 8
34475 vann 4
34476 vanor 3
34477 vansinne 3
34478 vansinnig 1
34479 vansinnigheter 1
34480 vansklig 1
34481 vanskliga 2
34482 vapen 23
34483 vapendragaren 1
34484 vapenhandeln 2
34485 vapenhandlare 1
34486 vapenindustrin 1
34487 vapenolja 1
34488 vapenrocken 1
34489 vapenvila 2
34490 vapenvilan 1
34491 vapnen 3
34492 var 1362
34493 vara 1198
34494 varade 3
34495 varaktig 10
34496 varaktiga 4
34497 varaktigt 4
34498 varan 3
34499 varandra 88
34500 varandras 3
34501 varann 1
34502 varannan 1
34503 varans 1
34504 varat 3
34505 varav 10
34506 varböld 2
34507 vardag 2
34508 vardagar 1
34509 vardagen 3
34510 vardagliga 5
34511 vardagligt 3
34512 vardags 1
34513 vardagsfraser 1
34514 vardagskriminaliteten 1
34515 vardagslag 1
34516 vardagsmat 1
34517 vardagspolitiken 1
34518 vardagsrum 1
34519 vardagsrummet 8
34520 vardagsrutin 1
34521 vardande 1
34522 vardera 1
34523 vare 100
34524 varefter 6
34525 varelse 5
34526 varelsen 1
34527 varelser 4
34528 varelserna 1
34529 varenda 16
34530 varför 121
34531 varg 1
34532 vargar 1
34533 vargarna 2
34534 varhelst 3
34535 vari 2
34536 variabel 2
34537 variabler 2
34538 variant 1
34539 varianter 1
34540 varierade 1
34541 varierande 4
34542 varierar 5
34543 varierat 1
34544 varifrån 5
34545 varigenom 2
34546 varit 318
34547 varje 288
34548 varken 47
34549 varm 4
34550 varma 9
34551 varmaste 1
34552 varmblodiga 1
34553 varmed 1
34554 varmt 31
34555 varmvattenberedaren 1
34556 varna 7
34557 varnade 2
34558 varnades 1
34559 varnagel 1
34560 varnande 1
34561 varnar 4
34562 varnat 2
34563 varning 14
34564 varningar 1
34565 varningarna 1
34566 varningen 1
34567 varningens 1
34568 varningssignal 1
34569 varningssystemet 1
34570 varor 21
34571 varorna 3
34572 varors 2
34573 varpbomtrålare 1
34574 varpå 4
34575 vars 88
34576 varsamma 1
34577 varse 1
34578 varsel 3
34579 varslar 1
34580 varstans 1
34581 varsågod 1
34582 vart 25
34583 vartannat 4
34584 vartenda 2
34585 varv 2
34586 varvid 12
34587 varvsindustrin 2
34588 varvsstöd 2
34589 vaska 1
34590 vassa 1
34591 vatten 129
34592 vatten- 1
34593 vattenanvändarna 4
34594 vattenanvändning 4
34595 vattenanvändningen 1
34596 vattenavgifter 3
34597 vattenbrist 6
34598 vattenbruk 5
34599 vattenbruket 2
34600 vattenbrukets 1
34601 vattenbruksanläggningar 1
34602 vattenbruksindustrin 2
34603 vattenbruksnäringen 1
34604 vattenbrukssektorn 4
34605 vattenbrukssystem 1
34606 vattenbrukssystemen 1
34607 vattenbyggnadsarbeten 1
34608 vattendammar 1
34609 vattendelare 2
34610 vattendirektiv 1
34611 vattendirektivet 2
34612 vattendistributionen 1
34613 vattendrag 5
34614 vattendragen 2
34615 vattendunkar 1
34616 vattenekosystem 1
34617 vattenextraktion 1
34618 vattenflöde 1
34619 vattenfrågan 1
34620 vattenfylld 1
34621 vattenfördelningen 1
34622 vattenföroreningar 1
34623 vattenförråden 1
34624 vattenförsämring 2
34625 vattenförsörjning 1
34626 vattenförsörjningen 1
34627 vattenförvaltning 1
34628 vattenförvaltningen 1
34629 vattengränser 1
34630 vattenhushållning 2
34631 vattenindikatorerna 1
34632 vattenkatastrof 1
34633 vattenkostnaden 1
34634 vattenkostnaderna 1
34635 vattenkraftsprojekt 1
34636 vattenkrig 1
34637 vattenkvalitet 6
34638 vattenkvaliteten 5
34639 vattenkvalitetområden 1
34640 vattenkällorna 1
34641 vattenlagstiftning 1
34642 vattenlagstiftningen 1
34643 vattenleverantörerna 1
34644 vattenmiljö 1
34645 vattenmiljön 6
34646 vattenmyndigheter 1
34647 vattenmyndigheterna 1
34648 vattenmängden 1
34649 vattenmätare 1
34650 vattennyttjande 1
34651 vattennät 1
34652 vattenområde 1
34653 vattenområden 3
34654 vattenområdet 2
34655 vattenpolitik 8
34656 vattenpolitiken 11
34657 vattenpolitikens 6
34658 vattenpriser 1
34659 vattenprispolitiken 1
34660 vattenproblematiken 1
34661 vattenproblemen 1
34662 vattenramdirektivet 1
34663 vattenramdirektivets 1
34664 vattenrening 1
34665 vattenreningsanläggningar 1
34666 vattenreningsutrustning 1
34667 vattenreserver 2
34668 vattenreserverna 2
34669 vattenreservernas 1
34670 vattenresurser 6
34671 vattenresurserna 12
34672 vattensaneringen 1
34673 vattensituation 1
34674 vattenskydd 1
34675 vattenskyddet 2
34676 vattenskyddslagstiftning 1
34677 vattenslöseri 1
34678 vattensystem 2
34679 vattensystemen 1
34680 vattensystemet 2
34681 vattentermer 1
34682 vattenterritorium 1
34683 vattentillgångar 1
34684 vattentillgången 1
34685 vattenutnyttjande 6
34686 vattenväg 2
34687 vattenvägar 8
34688 vattenvården 1
34689 vattenöverflöd 1
34690 vattnade 1
34691 vattnas 1
34692 vattnen 1
34693 vattnet 67
34694 vattnets 3
34695 veck 1
34696 vecka 26
34697 veckan 44
34698 veckans 1
34699 veckas 1
34700 veckobesök 1
34701 veckor 38
34702 veckorna 17
34703 veckoslut 1
34704 veckosluten 1
34705 veckotidningar 1
34706 ved 3
34707 vederbörande 2
34708 vederbörandes 1
34709 vederbörlig 10
34710 vederbörliga 2
34711 vederbörligen 4
34712 vederbörligt 3
34713 vedergällningsaktion 1
34714 vederkvickande 1
34715 vederlägger 1
34716 vedermödor 1
34717 vedertagna 1
34718 vedervärdiga 1
34719 vek 3
34720 vekhet 3
34721 vekheten 1
34722 velat 21
34723 vem 63
34724 vems 2
34725 venakulära 1
34726 venetiansk 1
34727 ventileras 1
34728 ventures 1
34729 veranda 1
34730 verandan 2
34731 verbala 1
34732 verifiable 1
34733 verifierar 1
34734 verifierbara 1
34735 verk 13
34736 verka 25
34737 verkade 32
34738 verkan 9
34739 verkar 114
34740 verkat 4
34741 verket 78
34742 verkets 2
34743 verklig 62
34744 verkliga 73
34745 verklige 2
34746 verkligen 354
34747 verklighet 29
34748 verkligheten 48
34749 verkligheterna 1
34750 verklighetsfrämmande 1
34751 verkligt 52
34752 verkningar 1
34753 verkningsfulla 1
34754 verkningsfullt 4
34755 verkningslösa 2
34756 verkningslöst 2
34757 verksam 2
34758 verksamhet 96
34759 verksamheten 25
34760 verksamheter 11
34761 verksamheterna 2
34762 verksamhets 1
34763 verksamhetsavbrottet 1
34764 verksamhetsbas 1
34765 verksamhetsbudgetering 1
34766 verksamhetsgrenar 2
34767 verksamhetsmiljön 1
34768 verksamhetsområde 5
34769 verksamhetsprogram 1
34770 verksamhetstiden 1
34771 verksamhetstillväxt 1
34772 verksamhetsutveckling 1
34773 verksamhetsutövare 2
34774 verksamhetsutövarna 1
34775 verksamhetsutövarnas 1
34776 verksamhetsår 1
34777 verksamma 9
34778 verksamt 2
34779 verkstad 1
34780 verkstadsindustrin 1
34781 verkställa 7
34782 verkställande 9
34783 verkställandet 6
34784 verkställare 1
34785 verkställas 4
34786 verkställdes 1
34787 verkställer 3
34788 verkställighet 3
34789 verkställigheten 5
34790 verkställighetssynpunkt 1
34791 verkställs 2
34792 verkställts 1
34793 verktyg 18
34794 verktygen 1
34795 verktygsfält 1
34796 verktygsfältet 1
34797 verktygsstålstillverkarna 1
34798 vermouths 1
34799 versa 1
34800 versaler 3
34801 version 10
34802 versionen 16
34803 versioner 2
34804 versionsnumret 1
34805 vertikal 2
34806 vertikala 4
34807 vet 377
34808 veta 92
34809 vetat 2
34810 vetenskap 18
34811 vetenskapen 10
34812 vetenskapens 4
34813 vetenskaplig 20
34814 vetenskapliga 53
34815 vetenskapligt 8
34816 vetenskapsmän 11
34817 vetenskapsmännen 8
34818 vetenskapsmännens 1
34819 veteran- 1
34820 veteranbilar 6
34821 veteranbilarna 1
34822 veterinärer 1
34823 veterinärfrågor 1
34824 veterinärpersonal 1
34825 veterligen 1
34826 veto 6
34827 vetorätt 3
34828 vetoröster 1
34829 vetskap 3
34830 vetskapen 3
34831 vette 1
34832 vetter 3
34833 vettet 1
34834 vettig 5
34835 vettiga 1
34836 vettigt 5
34837 vettlös 1
34838 vettvilling 1
34839 vevade 1
34840 vi 4681
34841 via 58
34842 vibrerande 1
34843 vice 34
34844 vicelehendakari 1
34845 vicepresident 1
34846 vickade 1
34847 vid 652
34848 vida 9
34849 vidare 108
34850 vidarebefordra 5
34851 vidarebefordrar 1
34852 vidarebefordras 2
34853 vidarebefordrats 1
34854 vidarebehandlas 1
34855 vidareutbildning 1
34856 vidareutveckla 2
34857 vidareutvecklas 1
34858 vidareutvecklat 1
34859 vidareutveckling 1
34860 vidareutvecklingen 1
34861 vidaste 2
34862 vidbrättade 1
34863 vidd 2
34864 vidden 5
34865 video 1
34866 videoförhör 1
34867 videokonferenser 4
34868 vidga 2
34869 vidgades 2
34870 vidgas 1
34871 vidgå 1
34872 vidhålla 1
34873 vidhåller 4
34874 vidhållit 1
34875 vidhålls 1
34876 vidhöll 1
34877 vidmakthålla 3
34878 vidmakthållas 1
34879 vidmakthålls 1
34880 vidriga 1
34881 vidröras 1
34882 vidrörd 1
34883 vidrörde 1
34884 vidskeplighet 1
34885 vidsträckt 1
34886 vidsynta 1
34887 vidta 94
34888 vidtaga 1
34889 vidtagit 10
34890 vidtagits 6
34891 vidtagna 4
34892 vidtalat 1
34893 vidtar 17
34894 vidtas 36
34895 vidtog 1
34896 vidtogs 5
34897 vidögd 1
34898 vifta 1
34899 viftade 1
34900 viftades 1
34901 viftar 2
34902 vigt 1
34903 vigvattnet 1
34904 vigör 1
34905 vika 2
34906 vikarierna 1
34907 viker 2
34908 vikt 47
34909 vikt- 3
34910 vikten 24
34911 vikter 1
34912 viktförlust 1
34913 viktgränsen 2
34914 viktig 223
34915 viktiga 196
34916 viktigare 31
34917 viktigast 4
34918 viktigaste 124
34919 viktigt 401
34920 viktklasser 1
34921 viktorianerna 1
34922 vila 7
34923 vilade 3
34924 vilande 1
34925 vilar 19
34926 vilat 2
34927 vild 4
34928 vilda 14
34929 vildar 1
34930 vildars 1
34931 vildaste 2
34932 vildmark 1
34933 vildmarken 2
34934 vildmarkens 1
34935 vilja 502
34936 viljan 23
34937 viljans 1
34938 viljekraft 1
34939 viljemässigt 1
34940 viljestark 1
34941 viljestarka 1
34942 vilka 269
34943 vilkas 10
34944 vilken 228
34945 vilket 614
34946 vill 1498
34947 village 1
34948 ville 86
34949 villervalla 1
34950 villig 8
34951 villiga 2
34952 villighet 2
34953 villigt 2
34954 villkor 85
34955 villkorade 1
34956 villkorande 1
34957 villkorar 1
34958 villkorat 1
34959 villkoren 30
34960 villkoret 1
34961 villkorlig 1
34962 villkorliga 2
34963 villkorligt 2
34964 villkorsuttryck 2
34965 villor 2
34966 villovägar 1
34967 villrådighet 1
34968 vilse 2
34969 vilsekommet 1
34970 vilseleda 2
34971 vilseledande 3
34972 vilseletts 1
34973 vilt 3
34974 vin 14
34975 vinade 1
34976 vind 5
34977 vindar 2
34978 vinden 3
34979 vindfällen 1
34980 vindfällena 3
34981 vindlande 1
34982 vindruta 1
34983 vindskyffe 1
34984 vinet 4
34985 vingla 1
34986 vinkade 3
34987 vinkande 1
34988 vinkelräta 2
34989 vinklade 1
34990 vinklar 2
34991 vinkling 1
34992 vinna 11
34993 vinnande 1
34994 vinnare 1
34995 vinnarna 1
34996 vinnas 1
34997 vinner 4
34998 vinning 1
34999 vinodlingar 1
35000 vinodlingen 1
35001 vinproduktionen 1
35002 vinsektorn 1
35003 vinst 11
35004 vinsten 3
35005 vinster 18
35006 vinsterna 4
35007 vinstinriktade 2
35008 vinstintresse 2
35009 vinstintresset 2
35010 vinstjakt 1
35011 vinstmarginaler 1
35012 vinstsvag 1
35013 vinsttänkande 1
35014 vint 1
35015 vinter 1
35016 vintereftermiddag 1
35017 vintern 3
35018 vintertid 1
35019 vinthunds 1
35020 vinylfodral 1
35021 violer 2
35022 vippade 1
35023 vippen 1
35024 vira 1
35025 virka 1
35026 virkesförsäljning 1
35027 virkeslager 1
35028 virkeslagren 1
35029 virrigt 1
35030 virrvarr 1
35031 virtuellt 2
35032 virus 4
35033 virusbärare 1
35034 viruset 8
35035 virussjukdom 2
35036 virveln 2
35037 virvelvind 1
35038 virvlade 2
35039 virvlande 1
35040 vis 30
35041 visa 101
35042 visade 32
35043 visades 1
35044 visar 154
35045 visare 1
35046 visas 28
35047 visat 79
35048 visats 3
35049 visavi 2
35050 visdom 1
35051 vise 1
35052 visering 1
35053 viseringar 1
35054 viserings- 1
35055 vises 1
35056 viset 11
35057 vishet 2
35058 vishetens 1
35059 vision 18
35060 visionen 3
35061 visioner 9
35062 visiteras 1
35063 viskade 2
35064 viskades 1
35065 visningsformat 1
35066 vispgrädde 1
35067 viss 108
35068 vissa 381
35069 visselpipa 1
35070 visselpipan 1
35071 visserligen 31
35072 visshet 3
35073 vissheten 1
35074 visslade 1
35075 visslande 1
35076 visst 32
35077 visste 50
35078 vistades 1
35079 vistas 4
35080 vistats 1
35081 vistelse 1
35082 vistelseort 1
35083 visualisera 1
35084 visuella 2
35085 visum 1
35086 vit 21
35087 vita 40
35088 vital 2
35089 vitala 3
35090 vitalisera 1
35091 vitaliseras 1
35092 vitalitet 1
35093 vitaliteten 1
35094 vitas 1
35095 vitaste 1
35096 vitblonda 1
35097 vitblänkande 1
35098 vitbok 34
35099 vitboken 44
35100 vitbokens 2
35101 vitbokssyndromet 1
35102 vitböcker 1
35103 vitböckerna 1
35104 vitglöd 1
35105 vitkalkade 1
35106 vitrinskåp 1
35107 vits 1
35108 vitt 15
35109 vittgående 1
35110 vittna 3
35111 vittnade 1
35112 vittnar 6
35113 vittnat 1
35114 vittne 3
35115 vittnen 1
35116 vittnesbördet 1
35117 vittnesförhör 1
35118 vittnet 1
35119 vittomfattande 4
35120 vittrande 1
35121 vittrar 1
35122 vitögat 1
35123 vivendi 2
35124 vokabulär 3
35125 volet 2
35126 voluntarism 2
35127 voluntaristiska 4
35128 volym 1
35129 volymen 2
35130 volymer 1
35131 von 23
35132 vore 82
35133 votering 1
35134 voteringssystemet 2
35135 votre 1
35136 votum 1
35137 vrak 6
35138 vrakdelarna 1
35139 vraket 3
35140 vrakets 1
35141 vrakgods 1
35142 vred 1
35143 vrede 3
35144 vreden 1
35145 vredgat 1
35146 vredgats 1
35147 vrida 3
35148 vrider 1
35149 vrist 1
35150 vrister 1
35151 vristerna 1
35152 vräkte 1
35153 vräkts 2
35154 vrålade 2
35155 vrålande 1
35156 vulkanen 1
35157 vunnen 1
35158 vunnet 2
35159 vunnit 9
35160 vuxit 3
35161 vuxna 6
35162 vy 1
35163 vyer 5
35164 vykort 1
35165 vyn 2
35166 väcka 9
35167 väckarklocka 2
35168 väcker 11
35169 väcks 2
35170 väckt 4
35171 väckte 5
35172 väcktes 4
35173 väckts 2
35174 väder 2
35175 väderkvarnar 1
35176 väders 1
35177 väderstreck 2
35178 vädja 6
35179 vädjan 9
35180 vädjanden 4
35181 vädjar 12
35182 vädjat 1
35183 vädret 4
35184 väg 121
35185 väg- 1
35186 väga 7
35187 vägar 29
35188 vägarna 9
35189 vägas 2
35190 vägbyggnad 1
35191 vägde 1
35192 vägen 71
35193 väger 4
35194 vägg 4
35195 väggar 2
35196 väggarna 9
35197 väggen 7
35198 vägkontroller 4
35199 vägkontrollerna 1
35200 vägleda 1
35201 vägledande 8
35202 vägledning 2
35203 väglett 3
35204 vägmärken 1
35205 vägnar 42
35206 vägnät 1
35207 vägra 10
35208 vägrade 6
35209 vägran 11
35210 vägrar 13
35211 vägras 1
35212 vägrat 6
35213 vägröjare 1
35214 vägskäl 1
35215 vägskälet 1
35216 vägsträckan 1
35217 vägsäkerhetens 1
35218 vägtrafikanter 1
35219 vägtrafikants 1
35220 vägtrafiken 1
35221 vägtrafiksäkerheten 1
35222 vägtransporter 1
35223 väktare 6
35224 väl 182
35225 välbalanserad 2
35226 välbalanserade 2
35227 välbefinnande 3
35228 välbehövligt 1
35229 välbekant 2
35230 välbekanta 1
35231 välbeställda 1
35232 väldig 8
35233 väldiga 6
35234 väldigt 69
35235 välformade 1
35236 välformat 1
35237 välfunna 1
35238 välfärd 14
35239 välfärden 4
35240 välfärdsmässiga 1
35241 välfärdsmålen 1
35242 välfärdsnivån 1
35243 välfärdspolitiken 1
35244 välfärdssamhälle 1
35245 välfärdsskillnader 1
35246 välfärdsstaten 3
35247 välfärdsvinster 1
35248 välförvaltad 1
35249 välgrundad 2
35250 välgrundade 1
35251 välgång 1
35252 välgörande 3
35253 välgörenhet 1
35254 välinformerad 1
35255 välinformerade 1
35256 välja 48
35257 väljarbastioner 1
35258 väljare 9
35259 väljarkåren 2
35260 väljarna 9
35261 väljarnas 2
35262 väljas 3
35263 väljer 23
35264 väljs 4
35265 välklingande 1
35266 välkommen 9
35267 välkommet 11
35268 välkomna 39
35269 välkomnade 2
35270 välkomnande 1
35271 välkomnar 88
35272 välkomnas 6
35273 välkomnat 1
35274 välkomnats 1
35275 välkomsthälsning 1
35276 välkvalificerade 1
35277 välkända 6
35278 välkänt 5
35279 vällde 1
35280 väller 1
35281 välmenande 2
35282 välment 1
35283 välmenta 2
35284 välmotiverad 1
35285 välmående 7
35286 välsignad 1
35287 välsignade 1
35288 välsignelse 1
35289 välsignelser 1
35290 välskött 1
35291 välstrukturerad 1
35292 välstånd 22
35293 välståndet 1
35294 välståndets 1
35295 välståndsnivå 1
35296 välståndsutvecklingen 1
35297 välta 1
35298 vältalig 1
35299 vältaligt 2
35300 vältra 1
35301 välutbildad 2
35302 välutbildade 1
35303 välutvecklad 1
35304 välutvecklade 1
35305 välvde 1
35306 vämjelse 1
35307 vän 24
35308 vända 24
35309 vändas 1
35310 vände 24
35311 vänder 16
35312 vändning 5
35313 vändningen 2
35314 vändpunkt 10
35315 vänja 1
35316 vänlig 4
35317 vänliga 3
35318 vänligare 1
35319 vänligen 4
35320 vänlighet 1
35321 vänligt 3
35322 vänner 27
35323 vännerna 1
35324 vänners 1
35325 vänorter 1
35326 vänskap 6
35327 vänskapliga 1
35328 vänskapligt 1
35329 vänskapsband 1
35330 vänster 25
35331 vänsterbetänkande 1
35332 vänsterkritiker 1
35333 vänstern 16
35334 vänsterns 2
35335 vänsterregeringar 2
35336 vänsterregeringarna 1
35337 vänsterregeringens 1
35338 vänstra 5
35339 vänt 4
35340 vänta 45
35341 väntad 1
35342 väntade 19
35343 väntan 15
35344 väntar 47
35345 väntas 1
35346 väntat 13
35347 väntrummet 1
35348 vänts 1
35349 väpnad 2
35350 väpnade 12
35351 värd 13
35352 värda 8
35353 värde 34
35354 värdedata 1
35355 värdefull 8
35356 värdefulla 10
35357 värdefullt 5
35358 värdegemenskap 5
35359 värdegrund 1
35360 värdelös 2
35361 värdelösa 2
35362 värdemässigt 1
35363 värden 41
35364 värdena 9
35365 värdenamn 2
35366 värdepapper 6
35367 värdepappersfonder 1
35368 värdepappersfondernas 1
35369 värdepappersmarknaden 1
35370 värdepappersområdet 2
35371 värdera 2
35372 värderade 7
35373 värderar 2
35374 värderas 5
35375 värdering 3
35376 värderingar 36
35377 värderingarna 4
35378 värderingarnas 1
35379 värdestegring 1
35380 värdesystem 1
35381 värdesätta 1
35382 värdesätter 1
35383 värdet 14
35384 värdeökningen 1
35385 värdig 3
35386 värdighet 14
35387 värdigheten 2
35388 värdigt 4
35389 värdinna 1
35390 värdinnorna 1
35391 värdlandet 1
35392 värdmedlemsstatens 1
35393 värja 1
35394 värjer 1
35395 värkande 1
35396 värkar 1
35397 värkte 1
35398 värld 30
35399 världar 3
35400 världen 163
35401 världens 39
35402 världsbefolkningen 1
35403 världsbild 1
35404 världsdel 6
35405 världsdelar 2
35406 världsdelen 3
35407 världsekonomin 7
35408 världsfinansens 1
35409 världsfrågorna 1
35410 världsfrånvända 1
35411 världshandel 2
35412 världshandeln 3
35413 världshandelsförhandlingar 1
35414 världsklockan 1
35415 världskonferens 2
35416 världskrig 1
35417 världskriget 5
35418 världskrigets 3
35419 världsledande 1
35420 världsliga 1
35421 världsmakts 1
35422 världsmarknaden 5
35423 världsmarknaderna 1
35424 världsmarknadsorientering 1
35425 världsmarknadspriserna 1
35426 världsmedborgare 1
35427 världsmodell 1
35428 världsnivå 1
35429 världsomspännande 7
35430 världsordning 3
35431 världsordningen 2
35432 världsregering 1
35433 världsriken 1
35434 världssamfundet 7
35435 världssamfundets 1
35436 världsstandard 1
35437 världsstyre 1
35438 världsuppfattning 1
35439 världsvana 1
35440 världsvattenforum 1
35441 världsövergripande 1
35442 värmas 1
35443 värmde 3
35444 värmdes 1
35445 värme 3
35446 värmen 2
35447 värmepannan 1
35448 värmt 2
35449 värna 9
35450 värnar 6
35451 värre 16
35452 värst 3
35453 värsta 23
35454 värt 14
35455 värv 2
35456 värvas 1
35457 väsande 1
35458 väsen 3
35459 väsendet 1
35460 väsentlig 17
35461 väsentliga 19
35462 väsentligen 2
35463 väsentligheterna 1
35464 väsentligt 23
35465 väska 3
35466 väskan 2
35467 väskorna 1
35468 väss 1
35469 väst 3
35470 västafrika 1
35471 västafrikanska 1
35472 väster 2
35473 västerländsk 1
35474 västerländska 1
35475 västerlänning 1
35476 västern 1
35477 västerut 1
35478 västeuropeiska 1
35479 västkusten 1
35480 västliga 1
35481 västländerna 3
35482 västländernas 1
35483 västra 7
35484 västvärlden 2
35485 väv 1
35486 vävnad 3
35487 vävnaden 1
35488 vävnader 1
35489 vävt 1
35490 växa 11
35491 växande 16
35492 växandets 1
35493 växelkontor 1
35494 växelkursen 1
35495 växelkurser 1
35496 växelkurserna 1
35497 växelkurspolitiken 1
35498 växelkursutvecklingen 1
35499 växelspel 1
35500 växelverkan 2
35501 växer 18
35502 växla 2
35503 växlande 1
35504 växlar 2
35505 växlas 1
35506 växlat 2
35507 växling 1
35508 växlingarna 2
35509 växtarter 1
35510 växte 6
35511 växter 4
35512 växtfrämjande 1
35513 växthuseffekt 1
35514 växthuseffekten 5
35515 växthusgaser 4
35516 växthusgaserna 2
35517 växtliv 2
35518 växtskydd 2
35519 växtskyddsproblem 1
35520 våg 2
35521 våga 3
35522 vågade 4
35523 vågar 13
35524 vågat 3
35525 vågen 1
35526 vågiga 1
35527 vågigt 1
35528 våglängd 1
35529 vågor 2
35530 vågorna 1
35531 vågrät 2
35532 vågskålen 1
35533 våld 12
35534 våldet 13
35535 våldets 2
35536 våldsam 5
35537 våldsamhet 1
35538 våldsamma 6
35539 våldsamt 4
35540 våldsbenägen 1
35541 våldsdemonstrationer 1
35542 våldsdåd 1
35543 våldsdåden 1
35544 våldshandlingar 2
35545 våldskultur 1
35546 våldsuttryck 1
35547 våldta 1
35548 våldtagen 1
35549 våldtagits 1
35550 våldtas 2
35551 våldtogs 1
35552 våldtäkt 2
35553 våldtäkter 1
35554 våldtäkterna 1
35555 vållade 1
35556 vållar 3
35557 våning 2
35558 våningar 1
35559 våningen 3
35560 vår 526
35561 våra 485
35562 vård 3
35563 vårda 1
35564 vårdad 1
35565 vårdade 1
35566 vårdar 3
35567 vårdcentraler 1
35568 vården 1
35569 vårdslös 1
35570 vårdslöshet 2
35571 våren 3
35572 vårens 1
35573 vårljus 1
35574 vårt 312
35575 vårta 1
35576 våta 1
35577 våtare 1
35578 våtmarksområden 1
35579 våtområden 1
35580 vått 1
35581 vördnad 3
35582 vördnadsbjudande 1
35583 vördnadsvärda 1
35584 walesare 1
35585 walesiska 1
35586 wallonska 1
35587 webben 3
35588 webbläsare 4
35589 webbläsaren 3
35590 webbplats 2
35591 webbplatsen 2
35592 webbsida 5
35593 webbsidan 1
35594 webbsidans 1
35595 webbsidor 2
35596 webbsidorna 1
35597 weitergeführt 1
35598 welfare 1
35599 werden 1
35600 whisky 7
35601 winschen 1
35602 with 3
35603 within 1
35604 worst 1
35605 yawlen 1
35606 yen 1
35607 ylade 1
35608 ylle 1
35609 yllesjalar 1
35610 yngelperioder 1
35611 yngre 5
35612 yngsta 1
35613 ynkliga 1
35614 ynkligt 1
35615 yppas 1
35616 ypperligt 2
35617 yppig 1
35618 yr 1
35619 yrka 7
35620 yrkande 6
35621 yrkanden 2
35622 yrkandet 2
35623 yrkar 8
35624 yrkat 1
35625 yrken 4
35626 yrkes- 1
35627 yrkesaktivas 1
35628 yrkesarbetande 2
35629 yrkesetik 1
35630 yrkesfiskarna 3
35631 yrkesfiskarnas 2
35632 yrkesgrupper 3
35633 yrkesjurister 1
35634 yrkeskarriärer 1
35635 yrkeskunnande 1
35636 yrkeskvalifikationer 2
35637 yrkeslivet 4
35638 yrkeslivets 1
35639 yrkesman 1
35640 yrkesmässig 1
35641 yrkesmässiga 2
35642 yrkesmässigt 1
35643 yrkesområdet 1
35644 yrkesprofil 1
35645 yrkestrafik 1
35646 yrkesutbildning 10
35647 yrkesutbildningen 2
35648 yrkesutbildningsåtgärder 1
35649 yrkesval 1
35650 yrkesverksamheter 1
35651 yrkesverksamma 7
35652 yrsel 1
35653 yt- 2
35654 yta 7
35655 ytan 4
35656 ytlig 1
35657 ytliga 1
35658 ytlighet 1
35659 ytligt 1
35660 ytorna 1
35661 ytskeendet 1
35662 ytterdörren 4
35663 ytterkläder 1
35664 ytterligare 189
35665 ytterligheten 3
35666 ytterligheter 1
35667 ytterlighetsåtgärder 1
35668 ytterligt 3
35669 ytterområde 1
35670 ytterområden 2
35671 ytterskrovet 1
35672 ytterst 62
35673 yttersta 34
35674 yttertrappan 1
35675 yttervärlden 2
35676 yttra 11
35677 yttrande 42
35678 yttrandefrihet 3
35679 yttranden 5
35680 yttrandet 13
35681 yttrar 2
35682 yttrat 1
35683 yttrats 3
35684 yttre 27
35685 ytvatten 9
35686 ytvattenstatus 2
35687 ytvattnen 1
35688 ytvattnens 1
35689 ytvattnet 8
35690 yviga 1
35691 yxa 1
35692 zero 1
35693 zigenare 3
35694 zigenarflyktingar 1
35695 zigenarna 1
35696 zigenska 1
35697 zon 2
35698 zoner 1
35699 zoners 1
35700 zonindelningen 1
35701 zu 9
35702 § 1
35703 ­ 1
35704 ­företräds 1
35705 ­inom 1
35706 º 1
35707 ¿ 1
35708 Álvaro 2
35709 Äldre 1
35710 Ämnar 1
35711 Ämnet 1
35712 Än 10
35713 Ända 6
35714 Ändra 4
35715 Ändras 1
35716 Ändring 1
35717 Ändringar 1
35718 Ändringsförslag 35
35719 Ändringsförslagen 11
35720 Ändå 27
35721 Ännu 11
35722 Äntligen 4
35723 Är 79
35724 Ärade 33
35725 Ärendet 1
35726 Ärkebiskopen 3
35727 Ärret 2
35728 Ät 1
35729 Även 123
35730 Å 67
35731 Åh 1
35732 Åhå 1
35733 Åklagaren 1
35734 Ånyo 1
35735 År 13
35736 Året 1
35737 Årligen 1
35738 Årligt 1
35739 Åsikt 2
35740 Åt 1
35741 Åtagandet 1
35742 Åtal 1
35743 Återetableringslagen 1
35744 Återigen 2
35745 Återinrättandet 1
35746 Återspeglas 1
35747 Återstående 1
35748 Återstår 2
35749 Återupptagande 6
35750 Återvinningskraven 1
35751 Åtgärd 1
35752 Åtgärder 10
35753 Åtgärderna 2
35754 Åtgärdernas 1
35755 Åtkomst 2
35756 Åtminstone 2
35757 Åtta 1
35758 Émilie 1
35759 Ésclope 1
35760 Île-de-France 1
35761 ÖVP 9
35762 Ödeslärjunge 1
35763 Ödet 1
35764 Ögonblicket 3
35765 Ögonen 1
35766 Öh 1
35767 Ökad 1
35768 Ön 1
35769 Önskar 1
35770 Önskemålet 1
35771 Öppenhet 2
35772 Öppna 1
35773 Öppnande 1
35774 Öst- 1
35775 Österrike 99
35776 Österrikes 14
35777 Österrikiska 11
35778 Östersjöländerna 1
35779 Östersjön 5
35780 Östersjöområdet 1
35781 Östersjöregionens 1
35782 Östeuropa 18
35783 Östeuropas 1
35784 Östtimor 8
35785 Östturkestan 1
35786 Östtyskland 4
35787 Över 6
35788 Överallt 1
35789 Överfisket 1
35790 Övergrepp 1
35791 Övergreppen 1
35792 Överproduktionen 1
35793 Överst 1
35794 Överste 2
35795 Översvämningar 1
35796 Översvämningarna 1
35797 Överväger 1
35798 Övriga 2
35799 à 1
35800 äcklar 1
35801 ädelstenar 2
35802 ädelt 2
35803 ädla 1
35804 äga 71
35805 ägandeform 1
35806 ägandeförhållanden 2
35807 äganderätten 1
35808 ägandet 1
35809 ägaransvaret 1
35810 ägare 10
35811 ägaren 8
35812 ägares 1
35813 ägarna 2
35814 ägarnas 1
35815 ägas 1
35816 ägde 14
35817 äger 33
35818 ägg 2
35819 ägna 24
35820 ägnad 1
35821 ägnade 8
35822 ägnar 29
35823 ägnas 4
35824 ägnat 9
35825 ägnats 1
35826 ägodelar 3
35827 ägt 15
35828 äkta 9
35829 äktenskap 2
35830 äktenskapsmål 1
35831 äkthet 1
35832 äldre 46
35833 äldreomsorg 1
35834 äldreomsorgen 1
35835 äldres 4
35836 äldsta 4
35837 älg 2
35838 älska 6
35839 älskade 9
35840 älskar 7
35841 älskare 1
35842 älskat 1
35843 älskvärd 1
35844 älskvärda 2
35845 älskvärdhet 1
35846 älvar 1
35847 ämbete 6
35848 ämbetsmannalagen 1
35849 ämbetsmännen 1
35850 ämbetsrum 1
35851 ämna 1
35852 ämnade 3
35853 ämnar 9
35854 ämne 44
35855 ämnen 62
35856 ämnena 9
35857 ämnesområde 2
35858 ämnesområdena 1
35859 ämnesprioriteringarna 1
35860 ämnet 16
35861 ämnets 1
35862 än 628
35863 ända 26
35864 ändamål 12
35865 ändamålen 1
35866 ändamålet 12
35867 ändamålsenlig 5
35868 ändamålsenliga 5
35869 ändamålsenligheten 2
35870 ändamålsenligt 4
35871 ändarna 1
35872 ände 5
35873 änden 2
35874 ändlös 2
35875 ändlösa 5
35876 ändock 1
35877 ändpunkter 1
35878 ändra 88
35879 ändrad 3
35880 ändrade 7
35881 ändrades 1
35882 ändrar 12
35883 ändras 27
35884 ändrat 10
35885 ändrats 9
35886 ändring 61
35887 ändringar 69
35888 ändringarna 13
35889 ändringen 13
35890 ändringsakter 1
35891 ändringsdirektiv 1
35892 ändringsförlag 1
35893 ändringsförslag 436
35894 ändringsförslagen 81
35895 ändringsförslaget 21
35896 ändringsförslagets 1
35897 ändå 165
35898 ängarna 2
35899 ängel 1
35900 ängels 1
35901 ängen 1
35902 ängslan 2
35903 ängsliga 2
35904 ängsligt 4
35905 änka 1
35906 ännu 243
35907 äntligen 70
35908 äntrade 1
35909 äppel-pie 1
35910 är 8406
35911 ära 1
35912 ärade 116
35913 äran 11
35914 ärende 36
35915 ärenden 8
35916 ärendena 6
35917 ärendet 20
35918 ärendets 1
35919 ärkebiskopen 1
35920 ärkefiende 1
35921 ärlig 5
35922 ärliga 6
35923 ärlighet 1
35924 ärligt 11
35925 ärmarna 2
35926 ärmen 1
35927 äro 1
35928 ärofylld 1
35929 ärr 2
35930 ärrbildning 1
35931 ärret 1
35932 ärver 1
35933 ärvt 1
35934 ät 1
35935 äta 21
35936 ätas 1
35937 äter 7
35938 ätit 3
35939 ättning 1
35940 även 822
35941 äventyr 2
35942 äventyra 11
35943 äventyrades 1
35944 äventyrar 14
35945 äventyrare 1
35946 äventyras 5
35947 äventyret 1
35948 å 92
35949 åberopa 4
35950 åberopar 1
35951 åberopas 1
35952 åder 1
35953 ådra 1
35954 ådrog 1
35955 ådror 2
35956 ådrorna 1
35957 åh 1
35958 åhörare 1
35959 åhörarläktaren 3
35960 åhörarläktarna 1
35961 åhört 1
35962 åka 8
35963 åker 3
35964 åkerier 1
35965 åkern 1
35966 åklagare 20
35967 åklagaren 8
35968 åklagares 1
35969 åklagarmyndighet 9
35970 åklagarmyndigheten 4
35971 åklagarmyndigheter 1
35972 åklagarna 1
35973 åklagarämbete 1
35974 åkommor 1
35975 åkte 2
35976 ål 2
35977 ålagd 2
35978 ålagda 2
35979 ålagts 2
35980 ålder 17
35981 ålderdomen 2
35982 ålderdomlig 1
35983 ålderdomshem 2
35984 åldern 2
35985 ålders 1
35986 ålderspensionen 1
35987 ålderstigen 1
35988 ålderstigna 1
35989 åldersökning 1
35990 åldrade 1
35991 åldrande 5
35992 åldrandet 1
35993 åldras 1
35994 åldrats 1
35995 åldringar 1
35996 åligga 3
35997 åligger 7
35998 ålägga 5
35999 ålägganden 1
36000 åläggandet 1
36001 åläggas 1
36002 ålägger 6
36003 åläggs 1
36004 ån 1
36005 ångare 2
36006 ångat 1
36007 ångbåtar 1
36008 ånger 1
36009 ångestfyllda 1
36010 ångestfyllt 1
36011 ånglok 1
36012 ångorna 1
36013 ångpanna 1
36014 ångrade 1
36015 ångvälten 1
36016 ånyo 3
36017 år 588
36018 år- 1
36019 åra 1
36020 åratal 9
36021 åren 127
36022 årens 13
36023 året 90
36024 årets 7
36025 århundrade 8
36026 århundraden 4
36027 århundradet 14
36028 århundradets 1
36029 årlig 6
36030 årliga 35
36031 årligen 14
36032 årligt 2
36033 års 42
36034 årsbeloppet 1
36035 årsberättelser 1
36036 årsrapport 3
36037 årsrapporten 2
36038 årsrapporter 1
36039 årstiden 1
36040 årsungar 2
36041 årsvis 1
36042 årtal 1
36043 årtionde 1
36044 årtionden 4
36045 årtiondena 1
36046 årtiondet 1
36047 årtusende 2
36048 årtusendena 1
36049 årtusendeskiftet 1
36050 årtusendet 1
36051 årtusendets 1
36052 åsamkar 1
36053 åsamkas 1
36054 åsamkat 4
36055 åsatt 1
36056 åsidosatte 1
36057 åsidosattes 2
36058 åsidosätta 3
36059 åsidosättande 2
36060 åsidosätter 3
36061 åsikt 76
36062 åsikten 8
36063 åsikter 37
36064 åsikterna 9
36065 åsiktsförbrytelser 1
36066 åsiktsförklaring 1
36067 åsiktsskillnad 1
36068 åsiktsskillnader 2
36069 åsiktsutbyten 1
36070 åskådarbalkongen 1
36071 åskådare 3
36072 åskådaren 1
36073 åskådliggjordes 1
36074 åskådning 1
36075 åsna 1
36076 åsnejacka 1
36077 åsnor 2
36078 åsnorna 1
36079 åstad 1
36080 åstadkom 2
36081 åstadkomma 39
36082 åstadkommas 3
36083 åstadkommer 7
36084 åstadkommit 7
36085 åstadkommits 3
36086 åstadkoms 1
36087 åsyftade 5
36088 åsyftar 5
36089 åsyftas 4
36090 åsynen 1
36091 åt 301
36092 åta 6
36093 åtagande 28
36094 åtagande- 1
36095 åtaganden 40
36096 åtagandena 4
36097 åtagandet 6
36098 åtagandetakt 1
36099 åtagit 10
36100 åtal 8
36101 åtala 3
36102 åtalade 2
36103 åtalas 4
36104 åtalsfasen 1
36105 åtalspunkter 3
36106 åtalspunkterna 3
36107 åtanke 8
36108 åtar 5
36109 åter 64
36110 återanpassa 1
36111 återanpassning 2
36112 återanställningsprocesserna 1
36113 återanvända 3
36114 återanvändas 1
36115 återanvändbara 1
36116 återanvändning 9
36117 återanvändningen 1
36118 återanvändnings- 1
36119 återanvändningsbart 1
36120 återanvändningsnivåer 1
36121 återanvänt 1
36122 återbetala 2
36123 återbetalats 1
36124 återbetalning 2
36125 återerövra 1
36126 återerövrande 1
36127 återerövring 1
36128 återetableringslag 1
36129 återfaller 1
36130 återfick 1
36131 återfinnas 2
36132 återfinner 2
36133 återfinns 6
36134 återfunna 1
36135 återfunnen 1
36136 återfå 1
36137 återfår 1
36138 återföras 2
36139 återfördela 1
36140 återfördes 1
36141 återförena 2
36142 återförenat 1
36143 återförening 1
36144 återföringen 1
36145 återförs 1
36146 återförts 1
36147 återförvisa 1
36148 återförvisas 3
36149 återförvisning 1
36150 återförvisningen 1
36151 återförvärva 1
36152 återgav 2
36153 återgavs 2
36154 återge 8
36155 återger 2
36156 återges 2
36157 återgett 1
36158 återgick 1
36159 återgivande 1
36160 återgivning 1
36161 återgå 2
36162 återgång 1
36163 återgår 1
36164 återgått 1
36165 återhämta 2
36166 återhämtning 9
36167 återhämtningen 4
36168 återhämtningsnivåer 1
36169 återhämtningsprogram 1
36170 återhållen 1
36171 återhållsam 1
36172 återhållsamhet 1
36173 återhållsamma 4
36174 återigen 50
36175 återinför 2
36176 återinföra 2
36177 återinförande 1
36178 återinförs 1
36179 återinresa 1
36180 återintagande 1
36181 återintegrering 1
36182 återintegreringsprogram 1
36183 återkalla 2
36184 återkallad 1
36185 återknyta 2
36186 återkom 1
36187 återkomma 6
36188 återkommande 5
36189 återkommer 6
36190 återkommit 1
36191 återkomst 1
36192 återkomsten 1
36193 återkräva 2
36194 återkrävas 1
36195 återlämna 3
36196 återlösaren 1
36197 åternationalisera 3
36198 åternationaliseras 1
36199 åternationalisering 7
36200 åternationaliseringen 1
36201 återsamla 1
36202 återskapa 7
36203 återspegla 3
36204 återspeglade 1
36205 återspeglar 6
36206 återspeglas 4
36207 återspegling 1
36208 återstod 1
36209 återställa 25
36210 återställande 4
36211 återställandet 2
36212 återställas 1
36213 återställer 1
36214 återställs 1
36215 återstående 4
36216 återstår 28
36217 återsända 1
36218 återsänds 1
36219 återta 2
36220 återtagande 4
36221 återtagandet 3
36222 återtar 1
36223 återtas 1
36224 återtog 1
36225 återuppbygga 2
36226 återuppbyggandet 5
36227 återuppbyggnad 8
36228 återuppbyggnaden 12
36229 återuppbyggnader 1
36230 återuppbyggnadsarbete 1
36231 återuppbyggnadsarbetena 1
36232 återuppbyggnadsfas 1
36233 återuppbyggnadsorgan 1
36234 återuppbyggnadsprogram 2
36235 återuppbyggnadsprogrammet 1
36236 återuppbyggt 1
36237 återuppfinna 1
36238 återuppliva 1
36239 återupplivande 1
36240 återupplivandet 1
36241 återupprepa 1
36242 återupprepas 3
36243 återupprätta 13
36244 återupprättandet 1
36245 återupprättar 2
36246 återupprättas 2
36247 återuppstå 1
36248 återuppståndelse 1
36249 återuppstår 1
36250 återuppstått 1
36251 återuppta 4
36252 återupptagande 1
36253 återupptagandet 2
36254 återupptagen 5
36255 återupptagits 1
36256 återupptagna 2
36257 återupptar 3
36258 återupptas 3
36259 återupptogs 13
36260 återupptäcka 1
36261 återuppvaknandet 1
36262 återverkan 1
36263 återverkningar 1
36264 återvinna 16
36265 återvinnande 2
36266 återvinnas 7
36267 återvinner 3
36268 återvinning 22
36269 återvinningen 6
36270 återvinningsbart 1
36271 återvinningsföretag 1
36272 återvinningsgrad 1
36273 återvinningsindustrin 1
36274 återvinningskostnaderna 2
36275 återvinningskravet 1
36276 återvinningsmodell 1
36277 återvinningsmonopol 1
36278 återvinningsmål 2
36279 återvinningsmålet 1
36280 återvinningsprocessen 1
36281 återvinningssektor 1
36282 återvinningssektorn 1
36283 återvinningssystem 1
36284 återvinningsverksamheten 1
36285 återvinningsvänliga 1
36286 återvinns 2
36287 återvunna 1
36288 återvunnet 1
36289 återvända 7
36290 återvände 2
36291 återvänder 4
36292 återvändsgränd 2
36293 återvänt 3
36294 åtfölja 5
36295 åtföljande 4
36296 åtföljas 8
36297 åtföljde 1
36298 åtföljdes 1
36299 åtföljer 1
36300 åtföljs 6
36301 åtföljt 1
36302 åtföljts 1
36303 åtgärd 47
36304 åtgärda 2
36305 åtgärdar 2
36306 åtgärdas 5
36307 åtgärden 8
36308 åtgärdens 1
36309 åtgärder 447
36310 åtgärderna 37
36311 åtgärds 1
36312 åtgärdsgrupper 1
36313 åtgärdsgrupperna 1
36314 åtgärdslista 2
36315 åtgärdsområden 1
36316 åtgärdspaket 7
36317 åtgärdspaketet 1
36318 åtgärdsplan 4
36319 åtgärdsplanen 1
36320 åtgärdsplanerna 1
36321 åtgärdsprogram 9
36322 åtgärdsprogrammen 2
36323 åtgärdsprogrammet 1
36324 åtgärdspunkter 1
36325 åtgärdsrelaterade 1
36326 åthävor 1
36327 åtkomlig 1
36328 åtkomst 1
36329 åtlydd 1
36330 åtminstone 95
36331 åtnjuta 6
36332 åtnjutande 1
36333 åtnjuter 3
36334 åtnjöt 1
36335 åtog 3
36336 åtrådd 1
36337 åtrådde 2
36338 åtrår 1
36339 åtråvärdhet 1
36340 åtskilda 1
36341 åtskilja 1
36342 åtskillig 1
36343 åtskilliga 3
36344 åtskilligt 1
36345 åtskillnad 5
36346 åtstramning 4
36347 åtstramningar 2
36348 åtta 15
36349 åttasidiga 1
36350 åttatiden 1
36351 åttonde 2
36352 åvilar 3
36353 ö 6
36354 öar 2
36355 öarna 12
36356 öarnas 1
36357 öbo 1
36358 öbor 1
36359 öde 31
36360 ödelade 2
36361 ödelagd 1
36362 ödelagda 2
36363 ödelägga 1
36364 ödeläggande 1
36365 ödeläggelse 2
36366 ödeläggelsen 1
36367 ödeläggs 1
36368 ödemark 2
36369 ödemarken 1
36370 öden 1
36371 ödesbestämda 1
36372 ödesbestämt 1
36373 ödesdiger 2
36374 ödesdigert 2
36375 ödesdigra 5
36376 ödesgemenskap 3
36377 ödesmättade 1
36378 ödet 1
36379 ödslig 1
36380 öga 8
36381 ögat 4
36382 ögla 1
36383 ögon 62
36384 ögonblick 57
36385 ögonblicken 2
36386 ögonblicket 24
36387 ögonblickligen 1
36388 ögonbrynet 1
36389 ögonen 19
36390 ögonfärg 1
36391 ögonlocken 1
36392 ögontjänarna 1
36393 ögonvitor 1
36394 öka 99
36395 ökad 68
36396 ökade 27
36397 ökades 1
36398 ökande 14
36399 ökar 50
36400 ökas 7
36401 ökat 40
36402 öken 1
36403 ökenområden 1
36404 ökenområdet 1
36405 ökenspridningen 1
36406 ökenutbredning 2
36407 ökenutbredningen 1
36408 öknar 1
36409 öknen 1
36410 ökning 32
36411 ökningar 1
36412 ökningen 8
36413 ökningseffekt 1
36414 ökningsprincipen 1
36415 öl 6
36416 ölen 2
36417 ölflaskorna 1
36418 ölkrus 1
36419 ölsort 1
36420 öm 1
36421 ömma 1
36422 ömmande 1
36423 ömsesidig 10
36424 ömsesidiga 5
36425 ömsesidighet 1
36426 ömsesidigt 9
36427 ömtåliga 3
36428 ömtålighet 1
36429 ömänniskor 1
36430 ön 21
36431 öns 6
36432 önska 21
36433 önskad 3
36434 önskade 8
36435 önskan 36
36436 önskar 57
36437 önskas 1
36438 önskat 5
36439 önskelista 1
36440 önskelistan 1
36441 önskelistor 1
36442 önskemål 16
36443 önskemålen 2
36444 önsketänkandet 1
36445 önskning 1
36446 önskningar 6
36447 önskvärd 6
36448 önskvärda 3
36449 önskvärt 18
36450 öområden 2
36451 öområdena 1
36452 öppen 35
36453 öppenhet 90
36454 öppenheten 17
36455 öppenhetens 1
36456 öppenhets- 1
36457 öppenhetslag 1
36458 öppenhetslagstiftning 1
36459 öppensinnade 1
36460 öppet 37
36461 öppettider 1
36462 öppna 47
36463 öppnad 1
36464 öppnade 13
36465 öppnades 3
36466 öppnandet 1
36467 öppnar 20
36468 öppnare 3
36469 öppnas 8
36470 öppnat 2
36471 öppnats 2
36472 öppning 4
36473 öppningar 3
36474 öppningsanförande 1
36475 öppningsanförandet 1
36476 öppningserbjudande 1
36477 öppningshögtid 1
36478 öra 5
36479 örat 1
36480 öre 2
36481 öregion 1
36482 öregioner 5
36483 öregionerna 9
36484 örlogsmannen 1
36485 örngott 1
36486 örnnäsa 1
36487 öron 7
36488 öronbedövande 2
36489 öronen 3
36490 öronmärka 1
36491 öronmärkta 1
36492 öronsprängning 1
36493 ösa 1
36494 ösamhällen 1
36495 öst 4
36496 öst- 2
36497 östaterna 2
36498 östblocket 1
36499 öste 2
36500 öster 4
36501 österländska 1
36502 östern 2
36503 österrikare 3
36504 österrikarens 1
36505 österrikares 1
36506 österrikarna 5
36507 österrikisk 5
36508 österrikiska 56
36509 österrikiske 2
36510 österrikiskt 1
36511 österut 2
36512 östeuropeisk 1
36513 östeuropeiska 5
36514 östländerna 2
36515 östländernas 1
36516 östra 10
36517 östrepublikerna 1
36518 östutvidgningen 2
36519 öva 1
36520 övat 1
36521 över 714
36522 överallt 24
36523 överarmen 1
36524 överbefolkade 1
36525 överbefälhavare 1
36526 överbelasta 1
36527 överbelastad 3
36528 överbemanning 1
36529 överblick 1
36530 överblicka 1
36531 överblivna 1
36532 överbord 2
36533 överbringa 1
36534 överbrygga 4
36535 överbryggas 1
36536 överbud 4
36537 övercentralisering 1
36538 överdimensionerad 1
36539 överdrift 2
36540 överdrifter 1
36541 överdriva 1
36542 överdrivas 1
36543 överdriven 12
36544 överdriver 3
36545 överdrivet 8
36546 överdrivna 5
36547 överdåd 1
36548 överdådiga 1
36549 överens 108
36550 överenskommelse 38
36551 överenskommelsen 6
36552 överenskommelser 5
36553 överenskommelserna 1
36554 överenskommen 1
36555 överenskommet 2
36556 överenskommits 2
36557 överenskomna 5
36558 överensstämde 1
36559 överensstämma 6
36560 överensstämmande 3
36561 överensstämmelse 19
36562 överensstämmer 22
36563 överexploatering 1
36564 överfall 3
36565 överfallet 1
36566 överfarterna 1
36567 överfiske 2
36568 överfiskning 1
36569 överflyttas 1
36570 överflyttning 2
36571 överflödig 2
36572 överflödigt 3
36573 överfulla 1
36574 överföll 3
36575 överför 5
36576 överföra 9
36577 överförande 1
36578 överföras 6
36579 överförda 1
36580 överföring 20
36581 överföringar 2
36582 överföringarna 1
36583 överföringen 5
36584 överförs 6
36585 överförts 1
36586 övergav 1
36587 överge 4
36588 överger 6
36589 överges 6
36590 övergick 1
36591 övergiven 1
36592 övergivenhet 1
36593 övergivit 1
36594 övergivits 3
36595 övergivna 5
36596 övergrepp 2
36597 övergripande 32
36598 övergå 3
36599 övergång 6
36600 övergången 8
36601 övergångs- 1
36602 övergångsbestämmelser 3
36603 övergångsbestämmelserna 1
36604 övergångsfas 1
36605 övergångsperiod 6
36606 övergångsperioden 5
36607 övergångsperiodens 1
36608 övergångsperioder 1
36609 övergångssystemet 2
36610 övergångsår 1
36611 övergår 6
36612 övergått 1
36613 övergödd 1
36614 överhanden 1
36615 överhuvud 2
36616 överhuvudtaget 8
36617 överhängande 2
36618 överhöghet 3
36619 överilat 2
36620 överinseende 2
36621 överkastet 1
36622 överklaga 2
36623 överklagande 2
36624 överklagandeförfarande 1
36625 överklaganden 2
36626 överklagar 1
36627 överklagat 1
36628 överkomliga 3
36629 överkomligt 1
36630 överkomma 1
36631 överkommit 1
36632 överkommits 1
36633 överkompensation 1
36634 överkörd 1
36635 överlade 2
36636 överlagda 1
36637 överlagt 1
36638 överlappar 3
36639 överlappning 2
36640 överlappningar 1
36641 överledas 1
36642 överledning 1
36643 överledningar 1
36644 överledningarna 1
36645 överledningen 4
36646 överleva 11
36647 överlevandet 1
36648 överlevde 3
36649 överlever 3
36650 överlevnad 3
36651 överlevt 2
36652 överläggningar 7
36653 överläggningarna 2
36654 överlägsen 1
36655 överlägsenhet 2
36656 överlägsenheten 1
36657 överlämna 8
36658 överlämnad 1
36659 överlämnade 3
36660 överlämnades 4
36661 överlämnande 1
36662 överlämnandet 2
36663 överlämnar 15
36664 överlämnas 5
36665 överlämnat 4
36666 överlämnats 6
36667 överlåta 9
36668 överlåtandet 1
36669 överlåtas 1
36670 överlåtbara 4
36671 överlåtelse 1
36672 överlåtelser 1
36673 överlåter 2
36674 överlåtit 1
36675 överlåtits 1
36676 överlåts 2
36677 övermaskinist 1
36678 övermekaniserade 1
36679 övermodigt 1
36680 övermorgon 5
36681 övermänsklig 1
36682 övernationell 4
36683 övernationella 2
36684 övernitiska 1
36685 övernog 1
36686 överordnad 1
36687 överordnade 1
36688 överpriser 1
36689 överraskad 2
36690 överraskade 1
36691 överraskande 5
36692 överraskning 6
36693 överregionala 1
36694 överreglerande 1
36695 överreglerat 1
36696 överreglering 1
36697 överrock 2
36698 överrocken 2
36699 överrumplad 1
36700 överrumplat 1
36701 överräckande 1
36702 överrätten 1
36703 överrösta 1
36704 översatta 1
36705 översatte 1
36706 översattes 2
36707 översatts 1
36708 överseende 1
36709 översida 1
36710 översikt 6
36711 översikten 8
36712 översikter 1
36713 översiktsplan 1
36714 överskott 6
36715 överskottet 2
36716 överskottskapacitet 1
36717 överskridas 1
36718 överskrider 4
36719 överskridit 1
36720 överskridits 1
36721 överskrids 3
36722 överskriften 3
36723 överskugga 2
36724 överskuggar 1
36725 överskådlig 5
36726 överspänd 2
36727 överst 2
36728 översta 1
36729 överstat 1
36730 överstaten 1
36731 överstatliga 1
36732 överstatlighet 4
36733 överstatligt 1
36734 överste 1
36735 översteg 1
36736 överstiga 1
36737 överstiger 6
36738 överstigit 1
36739 överståndet 1
36740 överståndna 1
36741 översvämmade 2
36742 översvämmades 1
36743 översvämmas 1
36744 översvämning 2
36745 översvämningar 11
36746 översvämningarna 9
36747 översvämningsbistånd 1
36748 översvämningsproblem 1
36749 översyn 8
36750 översynen 3
36751 översänd 1
36752 översända 1
36753 översändes 1
36754 översänds 1
36755 översätta 2
36756 översättarhus 1
36757 översättas 1
36758 översättning 1
36759 översättningar 4
36760 översättningarna 3
36761 översättningen 5
36762 översättningsarbeten 1
36763 översättningsfelen 1
36764 översättningsmisstag 1
36765 översättningsproblem 2
36766 översättningsproblemet 1
36767 översättningstjänst 1
36768 översättningstjänsten 2
36769 översållad 1
36770 överta 8
36771 övertag 2
36772 övertagande 1
36773 övertaganden 1
36774 övertagits 1
36775 övertala 1
36776 övertalade 1
36777 övertar 1
36778 övertid 1
36779 övertog 2
36780 övertoner 1
36781 övertramp 2
36782 överträdde 1
36783 överträdelse 3
36784 överträdelser 15
36785 överträdelserna 1
36786 överträds 2
36787 överträffa 1
36788 överträffar 1
36789 övertyga 17
36790 övertygad 50
36791 övertygade 18
36792 övertygande 15
36793 övertygar 1
36794 övertygat 4
36795 övertygelse 16
36796 övertygelsen 3
36797 övertygelsers 1
36798 övertänkta 1
36799 övervaka 18
36800 övervakade 1
36801 övervakar 2
36802 övervakas 7
36803 övervakat 1
36804 övervakning 19
36805 övervakningen 6
36806 övervakningscentra 2
36807 övervakningscentrer 1
36808 övervakningscentrum 4
36809 övervakningsformer 1
36810 övervakningsinstans 1
36811 övervakningssystem 1
36812 överviktig 1
36813 övervinna 10
36814 övervinnas 1
36815 övervinner 1
36816 övervinns 1
36817 övervunnits 1
36818 överväga 37
36819 övervägande 7
36820 överväganden 10
36821 övervägas 2
36822 övervägd 1
36823 övervägda 1
36824 övervägde 1
36825 överväger 12
36826 övervägs 1
36827 övervägt 3
36828 överväldigades 1
36829 överväldigande 9
36830 övervältra 1
36831 övervåningen 3
36832 överösa 1
36833 övning 5
36834 övningarna 1
36835 övningsflygning 1
36836 övre 4
36837 övrig 6
36838 övriga 91
36839 övrigas 1
36840 övrigt 103
36841 – 196
